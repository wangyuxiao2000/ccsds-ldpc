/*************************************************************/
//function: CCSDS-(32768,16384)LDPC编码器
//Author  : WangYuxiao
//Email   : wyxee2000@163.com
//Data    : 2024.1.229
//Version : V 1.0
/*************************************************************/
`timescale 1 ns / 1 ps

module encoder_32768_16384 (clk,rst_n,s_axis_tdata,s_axis_tvalid,s_axis_tready,m_axis_tdata,m_axis_tvalid,m_axis_tlast,m_axis_tready);
/************************************************生成矩阵设置************************************************/
localparam n = 32768;
localparam k = 16384;
localparam sub_size = 2048;
localparam G1_1 = 2048'h41FF744E6C2C8EEBDFE751F0E48E3018B355CE9FF5510EA4F619A375595F770BFF956F34CE6B303AEFFCA0B08D2AE1125ABFA44018D13D74521EFAD5C68EE2F3E7F820C3468AB9FB497D65F92FF4F532CE2AD26D469E5A4571760FE3C79645551BF8DA62D93C9163F455BF9B989808D4D2C4B51DE3F345FCAAAD1687E2CE2C60D53C5A93878FC64B21345EB8099CA63E6E3C3E504C4C2F57D821B4249B5F8470264DB447FB3F32FF512E7714545976D398A9FDF9D17EB21BE86B939CB1BF4EDAAEE9439034250612EFE0010663E1B0B9411E77D39CCCF1526B1D92F1019257E73F1B04544856F5F56362B829E0B8BCD3670F53E30C61CF48FFB4126C8B8FFB4D;
localparam G1_2 = 2048'hE7BAA3CCDF32288BAC2BDD1EE2114FC6D62C232AD06546891C8F987F95E7BA045AABB78E709EF3A8959F66D7C4AF068A2309A9077BD5D949CB82DF239E3AE5824313B07AC16A7CAF4361CCAB6AD87F783E53B8398E60E228CBD8A1DB628D58C82D7A409C3CCC1FEF2364A9DEEA6B26DD435E17F7741512DD9664BAF7AFF65F54C7A92595D02DCEA10BFB28404818CE28E3F3BDDF90F3A58183C53E21D4336273DC55F9943BA9E16CDE9FE6478AD9E3B2C0D26678A1990DEE8C45F9E5BCA5DEF05F423225A91C91283904B5C80F226231C760DE45CF4DD62D2335850FBD7B2B1FB75C905ED55BB86C79E3761A8DC735D6702EABA857EADE389B948AD6CD2DDB3E;
localparam G1_3 = 2048'h40EDE5EB12B4A9B1D0A77D140AEAA4C52386684FEB5261D6417DBE852AD75DBA8F3365B45DBE710B8FDCB0E7A7828A56FC2DA64D723475E05B6C6D90DD99AE06296DEEFC4307010B4E6122080C56E00022C4BD1C2477982441876138E633B9326306DBCF66E0E3F1BFD0A79EC9297115B0F82736CD509A0215BA3C781FE941CA722973ACB6F5288BE2467E5509A797D422D6A40BAE54720CB5EAEA06B8EE63AD8D67836DD38DFB7A8E2CCDFDF2C9824E0AA1B4E1D9F6F65154B6781800DB4BC7B6825BA9A2DB32C1650A1EA1F955DFF578283334ADB55B6923B5C18D73CDA4B8A1FC3DCC94CE7B3E61032FDDF6C02F169FC8BAB92325ED07C5140858C6F7C58E;
localparam G1_4 = 2048'h5CE73FAAC97099B51674FCA9BED14999A7A32DD37D043D3F8930C727C5AA8B1F44423401597678E5B2F8773EF42A9D4C8F6A2A50E555B5CC8BD0D6F5A11E920BEEAD7761FF2FB8D7B598FFB017C38419A7CF6F6EFEC9E42951031811248C1F02845E0863834063DA9792A940CC6048491580FA7C127A6C79DE86D1AAB57EED3C52E1689B9F0CB0B92A06CD44671E3CB09F6143C6DD8B4F334A2A8102BE717550A7BB8873ECD93FA38DDB637E051632FAD254B617487165482F002FD3176505A1DB8A74516C43C93753ACCC83E2582795470C8651DA2134780E8AAEDA5796C4D535FE012443AC3313E9FA49F314C7C46B91DCC1444E63EB4C7E5F175DAB205848;
localparam G1_5 = 2048'h534ECB2A510BD2789C0A221912A8E33704A2453CAA39FC39CA2757A6DB12DB073838635748A0F0652FEC51B01A6CFAA6392748ADC58CABE566E7DE2F323FEE0984BC9FEE73C14A599D543B6A57F32CF8EEAA4CAD92444D0983EB73A53FADB6666A170D22CA94FE64D4704D09D2E50BC3D38014B9CF300A54090B2A9D9FA7031DD42BEFDE0B8C6A32699D1D03FB4A301E4B6C852037B3826DACBB30C059B8076A5F134B191EF6A3A6D3673EA5702BB96D66728CED3ECA5EC10FD4C45A8776907E7D0FBF0299ABDEEDA262DA423CFBC97B1116BCEC5B0F524D5DB5600682D9A2032E8975661518479461C096E53E6AC6CBA0D63CDE94298625123EA12D3FE8ECF9;
localparam G1_6 = 2048'h7F2D33D537B2C386AD3FF2724C5DB36B09C03C28110D10708C41D35FCED5B4DAB73EAAFDEEFB27EDAE24C0875DBCB1BD3B517F3C2FFD0EA530FCE5238EE1D41C4F6B51F260BD4ACDC5AF5D93D278A9262EB036E662ABF46E6F0DC9076A325F87AF30F0CC1081E532F303934E71EBA6B554E27CB3E2C1D14806E94D34D9D1B42E7A8EDC68958AB62256402D84ED9ADB01FDBD8D29723B4B6FE12EDEBB2BB1810072E399ADA0D693D03524FEE077CD7EC77DBCBA8DDA5CE37558EF5729AF45B176017C25532509DDAC09D4CFFD496D5681E9AC6F3D8D3A8EF44498D1311F72D234E7C6D80E7F7EDFBA5CE498216603584564A6304C44D9D582E93F6B4A21E079B6;
localparam G1_7 = 2048'hA2812E5D9C4F5D675E347B3673E7A5BE487C0DEBFBA9CE4642C26152AD7CE2FED2916AEBFD486D2616830EEE9A9E5297D642316DD113D0A75296BDE81E23EF80E37680B637377D7748699E61A7EF04F58E22CB05FAFB72047B28BF99E8E6A4E5490519C1F9377A6081BA1EB2CB22EC06D29117C8EA95DC5008F6C37F41742BC16CCBD5636E81975573D0C33394BC0645712FB1C45EF400B02B462754B2B5E3C1B88DFF8B12D54EF73CA04A72A631F14BC0229349C672F030C59B7A30A035FFA9ACF5F584FE581B14BADA95C76A926C8715B61543AAE1B2F495442C4910DCC2FE13A48CE4469F7FF2A82B3809FAFD892C46255F8ED6E28DD0E4F4459BC62974A9;
localparam G1_8 = 2048'h2B4953E5ABEB175F44CA105A7ADEAEEDF43205E880FC132C1B541D73031EAF3D5BAE844C942BA146FBC2007EA7D03D21A4966BF78AEBA6DEEE0C2DECE0717512CA7EC376AD9E20310A62322569EA2E88234F545DFCE48E1EDB7E7F9D91D42A32372B2460E359F929AAFD5CCB256DC4FE6A0D41D5BD982EC04AC2E5717507562E2431A60A417C907C76CBCD967D70A9B30A044DE529516E6169337BDE6E584F88EA7ED5600393C0AD8CB9B016C16725AFA953F79783C47D3FF5044F52426E15AEBDBBAA33968C92049F78C909AE12D0C0BDC408301B60D6F1DA7BAE52452CD14357B53405CA591643B5BB7BDA2C319BD2AD69F76D78B8F93224392B5B1B8CCBAA;
localparam G2_1 = 2048'h5E9F8A36D54BF542282BBB890E99A67F313908AFB79F032F76D668744161AA6FA337D66FF8C5B6A739963831AD6A403C90D493308AF92B498E35948C6442FB787ACAF6D647719B2B8065437452BE7FE80C38BCF582819324CA59FDA04C5FD75D0B4AF19333483FC3E0F494F23F48107D77D0C84346BDB9CC4885D67B618D2A1181DAC5F8A62478A1367219B78DF044F8F4205E172E238D24DDEF095A4BA5A2E98620D0CAE04BA3070BCD2807ADEF51D6A6A36B85F9168C504617B27E055726F8330E64288CB632004E8F4805DCE49FFABA18FC9B4B905A41331ADCB31A08DE927A42EF4E1D41629E6200081C332DDAA1A9BB0AA41235DC75BE2B37A2FCF86512;
localparam G2_2 = 2048'h67688A4C1885A9AC447B90B905177539C45283CC12C65E030F08278DA67A80D3125E649085A2DCACBC6CD50AAAA4FD817F8EB9D2367F7B24A045DEA4D421F5311403B61EFEC93E8982FEE6FAADCABBF49BE6C33211EB8B87454F22BC6FBFC7E2A212BB072B032AD2886604A8AA1BBF838AA537E33626AB35B192664539E0749FF2D75E540FBEDF51D26F7AADE1C61838B27BE1174D9F997B37F45BAFE6A7E0C13E0CACFEB2271FE409030001CE926C88083BE86B71190F5C76C0AB544ACA7AA8957617AA9A25AC34089BC9B6C2955D76EB365C255789EB1C2CBE375732118FE793012413B8BD88AD3C40F12FB477D2CE0151A12C44B74D96F285BDBA24644A2D;
localparam G2_3 = 2048'h2E5CCA4FAC6E05C6F60F22DD7BF4ECFD738600B49D6E04C58B32472E86821C36D76830BBF7289864A87413957C99FDC33CB27322B415891C8EE37F2ADBFD7BE1742BAF90BC695684C2341F42783D63C231E5385397BA31A1EEDF51506CA2496C3159636AECEB12B2963E1A898F2DD5F7CECDBF9CF4A74C1DC34ACA81C2A15675056623C81693C719F5A581E7691B0AF4EE55F21E80337C5CBB9E5BC9718C16E1F2D21C2B1459D4E0BA4C3B58DA928A77D627F30ADB03372C60A40C46FA3EE2A17B7E08E4A1CEB38A71783FD68520A8DEADD59C71AB5866DBD89EEAA8FFEE2584A8293B3E838F5DF011A02EA602219096A637A40A3A52BA670F8CF52CEF8D1DD3;
localparam G2_4 = 2048'h2D5E2CD631CA6A7716D592C4ED79DC1AE5645E85E523705EEC3B5C5876F1E683E1EA4B3F7C3BFD2EDCDE26CA1000A2A4B9EBA72234D266E83DE349BFD4180C35308FD75168919CC484BF39F1F2073C0847370724ACF129A38C974362A06AD3B2757295EF9C9CD0601660B01975893B709A3193B8C5AA41271506224B860397086483A7A72871D608F912095B7708A6A43AAE6D46A29A32A9707E3764A31C37888B72B744D8C58F987B03F43E1AB2314B98363E81DE8B853E0FD3D1ACDC6C50C12D4E85F8687683362A16FAB585888CCA9142FFFE7ECB6A6888198D8624C594E4D5773A5E6EE00941622DCA192EFE3224C63D324C8D5E30A5DED6C8E7253CF4F0;
localparam G2_5 = 2048'hBACE39B799BE26B3AA88DEFD66F730FE5333314CB0DD2AAFD431CDEF4CD3104A82990F80703125C05D3EF807734E21999EC2588BEB68882FC1587C5E3E20C4514327671489714AE70220E16FE426F360E8BEFE11715D2687B0A4232AE728103BC00945CB9A4F000410C13525D00228904DD3E4237388DD3520E952158FD16625AB92BA1D19CAB202FCF6E46CFA7117F6EDDA508D21EE5913D2C9CBB85818E43247EF9608599D72401503AC1C912D8D883A76D7C19881FCA576F9A883A5061E91703E9893240249AF9236B4F5F0CC8243601CAB029A5B4B5AC20C3E6FCBFAEB1B5EBC065F48C72EA26DB805ACAE1070EF014BEF6E5168481F0D93E8B19B91E45C;
localparam G2_6 = 2048'h50ABCA6EC38986F5154435D24EDDC1C42162A6FD8004CE48F75EF46DFFAA48357B2FBF04C232DD1D94D8AA6CD477D7B38B3C2035C3E1240BEE678EC9FF216FFE0AF2B04C0B791FA9697D69D693F6FD269598209565A0C944B3813DCA80B6D1F6C936F594FBA2168706B5FD6E0C25FBD4A08A13B9F084DEC4D85AE66E17B7C714B2F57D6C0CAD1E366F5EDFE4F194F19CD4AC6F021FD7BBEB581E51C08E1686269E864D5E43879070F0AEFC87997B8D0F8418E1A388377A9FDDCE6C5DF864BCE214FA7084C097450F36F479C4E8D7ABEBAA1A4CEF7FBC32FD3B82310D55C5F8FFE6E7E2E48802DFEC4ACA4189F74BD74C373B889662812931A51392841B3B7109;
localparam G2_7 = 2048'h96F4161E8922BF7464D6C444F6E1A847AAA3ADA9DB8E89D0002D0F2FFD8F19A25C7A5D2E7D1AC1FE2493CFDFC5B5F25504E977ABAAC347E3A90853AEB8E0ABAB9607F9E0C2ABB73D8269F2D799E2DF98C5F3AA24B54F350F3935F7056469FC0C5140FC1D0093BF63F0B228E195C63E4B0925A9ED7635C14BCAB5CAE3F87E14F8C7A9591BFAF7DBCA13F0B3E158F71CFDD1D2B1B3E3DC43D118F9078535B389D7C3D7A98EEE583D0275B1F13AD3ACBAE657564452FA7FD093A05031720E17D0ABDEE26750F6EF6B5A7E467F6DCC9D53694B5710980481640854D5C2FCBDEB9C0BD24D1AF813116D7F43A1E5E26AA93A8C39CCC9404599EF04BEA49CB26F146039;
localparam G2_8 = 2048'h5B5DB2669B52E229F581E17DF01E63AC9250119F3E1AB74CD184F71FD4D3CDDBA6463953560988635C3D92DB08E3C7D5FD4AC8D79377F9EC2978008DC9B39683C9DF4B8F80324AAA93FD6794854D8C8AAA1D6F44E76C22ADE99A6B05541F23A2C0A4EEEE5D5E5A77F861070C719995725F9F512E82239672B73FE341788DBC43D2ADCAD5663315F001AAAB6B0223B5D38800BC5B84612A8C7363EB698075E78EA2AECFB9EA6F39376F3A84779DF1CD26206829D29F933AE96F4C58772291ADD4EB4AFCD2200997DF6E2756FD55D6880662ACFF4EEA2E2C109650305D2D77CC6AF698FD00BB4583216DB2BB7B862C46E63E0F33E475653B41556DE01A3ADA5AC5;
localparam G3_1 = 2048'h9D61E99E90B4A655DBE628512D71163B0D55CF890F0883DE290FE852765426984817BB000E424B30C9AC8AF36E7D02FE13E97569DC6272D7BC1808F64A4E5D82C68FD8049C568AE78858535E1610043E22185AC42F851E96D7D827B41DADF250B2CC8065ED363D4B79CACE3740AE5D78748A056BFA5D82CB541806004505222E34DC3DF2A931C78CF3E01E8B4239B2A777B5D316C3B7D1CD36A355F1B5809FF6F4179DF2BC04674A60678A15DB9C5E971FD3091FC723C6C6934F5A330F0942767462ED4299BAD314ABBF52C3DEA74ABA64FE0F35217D78DCB5E35F39CC7A90203D9EBB5657CF2B922481825892E1C0D0FA02776C57F681463588AE38B8F8C7E4;
localparam G3_2 = 2048'hEAD5D624BDC1767D9A76B395D9FF571424AA982D1B84D10B1FA210089DBDF4FA72BFE7E0DBB6E4FECDD177F39CBCC1E661334106F8832BAB53481612301AED316804D504C7FD323F90CEED68067519117BD902449DA9F18EF4C18629FADF1E8A2261E3E8B4ACBE5353B9F35F82B3DA3F5037B78031289D6EA0B1D28216A68FC0F5C4B8359D5B7B53B4D13BB2826F4C1AAE9AD15763580F86ACA3F8AF261C28632E5AE936979E0C5E7470B506FE72BEAB52EB9BAF209E17B76F3FADB409D8C26876F813B8C1E65B63B80E0DC1EB362AB68ECBEC1112616DA018DD648ED3339578EE9EDD010B98C598EE46F8294FB2D4194C847CA3668C4AD5C4F215CD528E7ABD;
localparam G3_3 = 2048'h8D99CA3AE5E78BE9BC8A4FE85A1F74BB26885B70C22197CB4B4975E38A7D35792FE89D822AB02D023CA2E4B3993CF4EEC735DD83BA840F781968D86FB40C97E8BA166E90EEC00D5C0165584A4A0BA2E011B7D6130FA9165D1AADE4B0A2051EA39BD32701D324E5DF9E4B139CA6748912F4723313502E1583F94184B6F5671670813C907BB87FE6057831AEF4BF8EA7C3DAF18DFBB14B85498616C8E9BB5DACA67A6B99827227D257C8A07978330AF16672F810827875C1FC16EB88CCEAE10F3E944EA299D57D6D339A75EABD0F63F611414C016FAFB43D9D8319E634BDFC2FCC68F667D003A81F68CE660C95DD4C655698A5C4C7EA2EFB225104851BE180E223;
localparam G3_4 = 2048'hF08980189A6EA5686BDCBB1DD7DDA79DF9D5A3E57DD1DB0D72E04CEDC96A1F536D096473D0F6F50EF026D0F945DF02B6E0CB8FA21497A0F300BC8E56C820230DBD59798B042594D6DDB54596C29FB8AC8ABBE97F2DB2575C3AFEA6DFBD52821A1F1BABACC65A67EA4D4F9985312D623D421819CE95E5AC52ABB1CEF1624FF062579AA42DF5FBA0524EB10829E3B1ABE19A8AADE7339CFB18A6F6A1F1F95FF0FD5E8BA08758AB6C5E2F59396C27826112942ABE831107A09C019875A9C736F174CF79876BC66123FA0BBCD12B690AFFCE6BAD86FC74732C71A128399280A19FA900873928605AB04A872C43307E8B6EE8B5A877C32FF940D4107CBB70B2A8E2F6;
localparam G3_5 = 2048'h2BEB5D055A4F4D2C7700CB1C4CF198063F5620D2FBE171D115228E7345CA518590D966EC97E8AF9F91CBAE57FD2A1FAEC8DF3B6B5EB209246BA063DDAEBF225C2AC19DD86B6CD26046BBE821A56ACCEA5F02EE7D99F741AA3BFD16F7143BE27343E4561901B6E35049EAE57D3088161A081AD7DD9D513D2F16162CE8508E3CC518D0406D5140B857B4E8AA32B91E8D7E2E81F367890339EA347F6A637B77FE205257DA53C3AA6790A030DB82A131CFCE7BBC2478746516A4F3AA3BA4F7EEF50B093D757BF3A906AE335B6A57AD393FE72D45D4E1399113EAA70916D0D18F69E1546DC660AC848F29DDF6E4C26B2370B88E8F16FC257DED35F084AB05D5715897;
localparam G3_6 = 2048'h29E88AAD50DD6E1643C4BB5B7659928FEA1F4D071ECA6FF18C33BB502E2930662F1A28B83FC99BA1475C40A028BE3FD9595DB4E128BACE3697D82E5FB74EF6F52E766071DFFDD617E7493D2E863ABA80C7B67C28402F5A4A5AFE349E66C1E4E2C03E62685AB692E7494CCAD1ED4436F99F14890EC1963085FF020BFC65099ACF664BA133A6029D981633D9AA2E593C8B0B96989A1F71AB9A04A12E58C73B5466470FFBC0ACC2BE4AA73FFE0EF76781B046EAFDDA61F8B87A6C2C988FB7334B0ECC0438A50BBFFB8DEEFBEE314F16262EB84DFBBD65DE19DA9163BDF97FE10BCC0B926812D9E81E03FC77DE38C9A6A079228B895B5CB65858D9ED1BA7CEA7AB1F;
localparam G3_7 = 2048'hEC9E78F6F3FF46589D589E93639B755C6C8B4236AF3D118A0E2D9E48B9FCE58F99B477277BC7A3848FC8F650C023FA93074C737CFC7EEB639A7DC8680F9E8FD14D74CA364A52947703DFB74E5C7354F2FCE7D3AA2DDCD71C720D94D855095D5963E8037AB2DE386CDC13B03B4341E5DCBBEF8D243CD54299B7D2CA76813663DB0A86A2371B3C9A6F8AAE57E5FCDE2FBFD8600944AA506A176194E10C3730DAE1A44C3979573E9BAD3D694ABD650788ED3BBAF0231FFB8A97003EC597F5BB39CB6FADB502C8370DBBD2873FF156859D591295B364FCEC40D2A1012E82940697EE78C4394297C4060798A9A94834C35A3B991A4A913BA1A28098DEBFD40FC00F37;
localparam G3_8 = 2048'h17112E14360FB3C7985E6AF149DFE4B2BF65C781F3DD99F8E8B95E7BD2156EDFAEDAE7ECB1FC1D4F2783B0EAFDE9CC7C54C165C176E1DDEEC61804E57778FE674DCF7B85BB81061C28BB692018205167305E7DEDDA36D70B39F7A48A45E57F7ACBE59F292E20C156E282F9C0E30D5CBFE071914C25F615A308FF4AD731777A7BA1C4D3E3EEF751118C7E15066033F58893EB04A26AB0FACCF2E778CD35EBC161DE0116759E956037A2A4ACB9DECAD6004C9AD4892E5FD3ECCB5D561B9D1BC953E8361E1197293A5AB030E0C513DA444B51AE022B999FA9B32A6CCE3F7BF364C7D2CA6049F2CB3863A627ECB2CE6DB3208AD18FC134D43430D782873B721047E2;
localparam G4_1 = 2048'hC2B13C6F23387B4B65F28DF95A3EED6A7A1C3C49B65F3E9034E7A2446B40F6718AC1AB61F8D8ECE26F95EA795074FA1F95C4E149D2F7A5CD3A93DA0ADFE14DD257990D7588B87135FDA1275C6F3390073C7971541574159F1EE057C8A0BA227A16A0A93BB0E0C72DB8E33FB57A572579E0202B8E3DCCF2E42D2FC1255741FC24AD34E5EDDFE570450B7CE25378A7B61B94C4B0BE16492502BC5751818A0D5C9BF3EBAF11C78F74CC96EE284F235501F47D16A953C61BDD144B7E63EB9B8D719285BCD2374761BC201660A075107060135093B119F23BEACACA54022787F9169853D5963003EC43962F29630685BF7A6C35E177432497C547D250546EAA18963D;
localparam G4_2 = 2048'h4448FE5866E0C3ED55882CE597E0DA26689C07BE2D18CB6DD0F82CB0866747825EA19E8201F4EBB3ADB40677AA7D4C7D981141472C2C5CA77FC3B907BA9DA86C3D25A69A32494689B9E009318D36222F152D1DBFC82E65F87EEF063F9E68701833B889695467F1DE0594F71FA7B87CBE76EFFFA75E89BF2A69D4853A376BF38015D21FCB0B865B5FF94E383B322752FCBA04734280078171A49AAB0A22D2627AE030BC40A73319F84ABE65510A043DDBB6078C84D1F97DF693A7E8D55347FE1D5BACCACAF8DEEB7310E90B3FD3326CD3E17739C08291F1936FCB5C6CC5E9538062A9CCD83840D7864E500F1C31D7773F78BBBD6CE790854FD0363194B7408CBE;
localparam G4_3 = 2048'h4A6A8AE2595611E479893BF12D0ECEE5213AC2D1655214C5991FFCA99454CB51B377EA6AA7EA26EA0AF1000719DF1664857F14B7FE458EDDEF8ED24A175175F58260BADB642BA2562033ED084709B962D1E779F0E30FA1ECABD6C5FCB017802939C3890A77D38802BA064FCF78FE0FBCC06ED46C0E84C616ED95921979D7BAA2AF3041D761D1F095C41C875DFB0281F6971BA49BD2734D23D8EA08F254733F4B4C81265B330F47E9453DDE36EBBAE1EE60C0B0B3C8E0AA36184DCF477DA56C1601761D140205A36C9BAF5A7B724504777BE9D120B61BB67E678558551067CD3B311360E57E57A39EBC526302EA7598ECA0A4B0EE51AF04B73221A4F851B2098C;
localparam G4_4 = 2048'h3DFC370C05AE61AD51BD39A33469A077583EC0EA5D62892F56979664806EA9E61A3A4EA6CDDD9C7234BB9752822C55E8B0AA2007A2283BD0C5DD8DE70DB2BF1BBBB954C981760C64824ADB174A49BA5B7DA3EDC604EC269FA311287E9387A9E0EF8E16526418EC84648C5A0B040343A88CB8BEFB0E57CF5E66DF980A348816D12CE1A07DFDAEB9CC5D73D5D81B0CA56A0BC6785729F9080F41BBE35984AC428B48E1E98DF95C6BE71CD6B1DCF0D9A4A6CF9D9E4FF9BB58EDE3E1BD9AC3CF5BE495D6B0AE03CCEEA2154D8E16A514F37E312161B8137DA9ABEBC775EFE3D97DE570E8CA2240E30CFA6C05ED36527D6A3F6DC5867BFFAFDE85D0FBD24DBA34D25C;
localparam G4_5 = 2048'h740C3028574B45ADACA9657FFBEBA5996EB4FFCA666C2AE8CC180594C1B7FCA36391F5D68DE5FD3103256D572473675EFE1EE5CEF6B34D89A2F63A2CC68A20CBD965536EE4A2C33E3875E1EE368CB8FE74D21FECDB79381748900ACBC604A66CD8E8AA4FDEEECFEBAE2D3F305E51C5ACD33BE501DAC20704F34EDBF503E620E65ABA3906D695144AACD1AF7A6E716AF631BA1B5CC156FFE88109BAD0E324135580F327FA0308E72E2A3CA77C8848317E83D59CBDC239BBB5760E21605F006D0E0DA0B964D13F4FCD3AA9632F9EB7F21300FE284AC248CF8ED6AE15D2F177A3B801A5C8E3FEF0D5CBBFEC1FDF2E3F35E9A653530721D46B0BE576DDCE2EB7B6CC;
localparam G4_6 = 2048'h770969E2078BB0D1EB605A46FD651FB9C8933129A7058946E88C48BAF86350EC0F413FDCD2B3A9875A57B920B69157715D8CA707D15496D9DD19FB6F9614678119B34E676C44485D4F84CA5D5F8AD864DE2956C104A791F4B8928051C465758CBFF358B39799D53221DB3ECD6059EDC6C2E785E98FFA5BEB282C1F0B209953ADEF4A9B8D3A68D1D8E20EDA29CB9F4521A646D1630060DF96967746C34ADF7D56AC172ADFD654B0C4FAA44FB5DD21175BF7AC05676F211233324358B9CDABC64995192FE6FCED61BA61A4438156BF5E33CF676174FA95F20F0927BA88338228099BFAC9BEA0C0F15CAFF72235C133E1974D180C6E8C7CA3D0A1BF772FB5530F6C;
localparam G4_7 = 2048'h11F5B2124E781BDFF110C1DD5D24BF6E7FDFFB361823A89589654518429D6E8D480C2C7401880620A03B8AE5F6DA4EDEA1D736FDE2FCF951B54344675037424AB0FD3C1E994C1E7701F3AD7E1121C6C730988C2E26E586F9AE6AD1180F31664F3991F95FB8C277FE4F1F7A3508ABA71F92553A6FDDFBC81A95C2C03BD725CAFBDBB524DD1FA2D33BA5C2A1EE4A73711604C24BFC76189C6F87FDDEADDBC41F83471116DD656AEC88425B9E26D49731D1A6A52CFE954B6FA08CA040FDF27518CBFEDB692173B017286870181E1709B72B335EE552A3A5AAD623A2250A658722C6A2A5001F1AFA7AC400AAD5B49E40D662326E232CF500AA9AC954BB2B99831967;
localparam G4_8 = 2048'hCEAC6F8A6D91F0E73962EC35A8A7235F6516502CB3C5FE0545865DCA4D611FBC225AC4344F4DF4402FB2A240633B48C51C9ADB284DF3A7DC701B733F151FC765E9D97C65C6EA96759D78981113F564D23900281932327CD7170E3DCF4D52D28ABC0F0ECF7980BEE4CD5DFFAA48A29C22FBE502B1149A15294AB91BB8F7E32B6566F9F1A87975132A9BD35F19621E55EDF4B00045C6E84FDB0B36B363687E42C0EF4179EBA8B372E8FF1DC59BA012CD4575EACE5934EAAC5EC90069EA19380A8434A8D125EDBD629EEA5A71169D31B93001571459CCD8E047690A09BDEF391341053DDB52A53DF7D3346A3124390AC602B21E821385ED9B6AD254941E3827F205;
localparam G5_1 = 2048'h8BA51C8707B4CF2F3CD5BC23F67A783DAB62EF89B9A92E270BE5879E585B38FAFEC62137F081A07071410A22099B34C4DF1E6E4B915C74632CB5CA25AACA5DD19F3E493631F7654C34AF6B6CF5B93CB1EF59006E19A1D149649634F53455F842C2BDAB2FE836E79B76EF51C5D820E9EDED70B36CA00131EB2E2836477B4B89A51B0E3AA87DFDD32EEBD7824B8D4C1498000055D03A0DF344396B20FF99F4737BE4F94D7387051735E9C446FA69B5C7CB12F539CD7069844E515FEB95B0DCD0CAEB388B8E9C141141640AA944C73A7A69D6CAB7DA65DBEA3938C3D715EE7A7CDB58FCAAE768CDD87DA2B94E875B6696BC714385A9DD0372E157B8BB194A9962A0;
localparam G5_2 = 2048'h8503BCBD2A7D626B421CCF47344A03C802C8E050C7D9E4852602B05F475F1EED68B664D268E797F8FDEBA238485C3E125CA2D60A352635ECCABD983A6472BAD8E5312E79BF66FE94EB3079268AB5DB9B8CA174A28A953548948022F2F4914E8623CB75B3F1D1F70858A0CB42F8B86EF41E10099F354BF70C2D3C77B016251561A05B3E3F29098400D9109576F745A26795BE9BB1226D529CD3C5627088F2E79662F12CCF097B3FD5C23C4D42D396811C96E4FDC13F42DDC1D7A706BD34D79EB38571A5F24CF08314457F324F4AB4B39558FF13A04CB8B519E10E72983AD501ED90B268BCB08AE90D5413D36CEF7B4520F1DD7B9B15B6F369D710BE482E81AB98;
localparam G5_3 = 2048'hC7DA20EB864E02E959D9FB734E98215E2C50C926FA20409BBC2E4EB8EF13CAE99EBFDE473C0444BE0AAABFCC3828B97398A58AD2911074C45B24FBC4AB907AA6103A2F497554D5F7AAE399228C802B11C56C311A00C184C138B0FCFE97A1C278C7F0CC6C8FA479A73D7C6407E3AA7EA017E5652358033F0224E3DB2FEA069AB51CBAEFEE7E241AD1ED3679894954F7C0A0240403EBB32DCFCAE043ED9DB067DB56637BB124CB4E2C556FAEE519745762914E200B0CB5F38E463869777D6200343DC5D1B62E69E64D47E3D695337FBE286B4A506EB180CD44D637945F945B84A3C32A4C31501268CB14369682F63CF2EF788B0FED62FB35B1F3B1E10C06F7481B;
localparam G5_4 = 2048'h711E28BBAF6916C647A269BA5A072439A32CD6C24316C790D81892AF4FBAD18C834371FBB6A0397A8A1B078FD170B7E0385C2AB7FC2EED86262D93CC1E022A8954D5D58276345C536977B4217ADBBA97DF6A229EF423DE152559F033ECE4EBF8E3F5A5599723ABDE5F5639A2DD3BBFE673D35F1E2CFD872CC1C01044883038AF738AB66D339BB8A6434333211422348E7C8D33EC6E27FE772274AB9C8BABFF3C4A66C3767DE20B26CE0F042160384939A963ECFD5F0648577D30C886C3B73665745BDEBDEC5C9ABFE862E3B11537D482B79DCF2FACF08153E8A8AB2EB7174FD6FA879B6453D563E50CC27D844AD8F5B445E1E113689FC7117F89B177A2C7E6FA;
localparam G5_5 = 2048'hAC383DDC30B5DD262D17A541B605C83FAF6F7BFAA942C23156AD2D09CF5C62AD04AAB88324D941C6A755FC5DED8A80CCC15B90C45C53CA04E6995A738393365C102C5315FD1CB46019374C4A75C12CC1C393BA42EAA24AAC61471AA3222EB3E1D261B32F8F60142E88C3E3C413F87236F6C154FC25F7F41F9B8BD2EC335352812C31CBF8E0D4CFD76AAF50916BF3101410C729743E91DB515226B34094EF48E8AD7317DEA62C72735098A2DCC967FC2FBFC0E2609E6602DC34BCC1C15AA110EB015D780EE742C096FBAD9D2F2A0F698307DCC40D0CFEADD0C0987C96B2759D4CBE7B3A9026D58836639973722D6CCF2B1F98856AC3A4660F2A00412E8BDF06D8;
localparam G5_6 = 2048'h8732121CF94EF78889F383001FB85BBFF5187869F8A6CCA88A7D9D420A468868D09ABDB940F58437863411617C9B7E7984DC064804F5B61D576EF4816ECC3A22F265E1B258A2F5C1BDA6CB6D7A3C7B6BDAF2E6285037C1AD284B5375F023A5175996A85A086D7192CE47A50851F0FB7E568235BC68A8E8B8FCCDD6A0429BBE072F97F4359AD826F014743E43324CF65D1C7A6CADF08359CFF70DE3DECEE87BB29A247B9D463679B4313C1953B2E1B596704A25A85D8C694DFC7C91D73482547460029042DC89252570309A923F4651679695AD17B533435A211A7C6F83BEE182768812C12E928A55008AB724629C7BF5EFC5D02CC3D885F30E69AD27F17B80D7;
localparam G5_7 = 2048'h0BF5736667A2A2FF17AB3FD0F4D4350B006B20770932BCD2C64A91CA1CC307D7EE3AF75CEBCF4709765E74E85FB724D7EC5283F79C1573EBE23F510B685B99294790D43E0D45AFC213FE1FCC6DC1C2A53E8129DEF24BE5C27E7072F5EA1DDCC2B2CAD1334902EE3B7B0A907955D2B836AB5BCBFD4E250BE9AA8A2E0F896B6EBEC32135B878830F3C24F202F9925FFE2B0D6977F7A8E2010D9B18CE3E632335B084E7E2DB40064FE74197D384A694CFA6A4D1D855C8AAE51F7511EA7F1AB1A8E67AE10C02FB5C8117B56822072147F2A3813CF759146DAC0EEB4D48430250BE158F511AFDBE6F8CDB87B56C84AFF752812A7CC18BF22146F2B3AD6910B919EBDD;
localparam G5_8 = 2048'h37DD07C903337789882AF8169E6B1FC9396ADF225929E11BA5088AD37F83574C6F6579475F5EFA303E45526780F59D433405CFBC5EA28DEDD0A46E65CC3EA56581AC24F1495082ABDD3D320F777EA66BF9B6000DC0CA9082DE0EF5A18B7F7E1F98C556E29FC9B32DE74C94938C2661134B5E9B158F77C4641D856B5AC1B91FA7371BCCF1B80858F190F49CE920841AEE5EEDF74943D1CA8B9672022198AD911E4627D374A047C12C196457E2574D45708EF8765FE0DE1C4B9C48E1040F43E44D8BC8962170EDF6154F7E412C959A083854D83AACEADCE8058C8276F747DB7C71D0CB7DCF4A3D37882985B0A3CAAB2576D7EE195AC4292596E1397E44E13D09BA;
localparam G6_1 = 2048'h4AE7D32CA99DD4A718EC7998C5CEA77F65784558D31796FB5523E806608214ECBEB7F984FF5F15B8273ACEC88361194DA2AC962E2779AB50242D05AD9737197534268C0BDBAF84D2B962A9FCFC2375FEA2068C94CB1DB52ADDA678CE7865059118E7C2A6F69D3C17ACF48EC0C33CB35D14F92E2F574EEEC15DD28CA6341369C4B236088E1F3438FAD737C27E354F672FE86951673C17F88E62697DAEC5A4FB103A18FC5937C53B29C62BA6A973639441972B0E29F0A02F618CCB752AD3B8A468E8BE28F370E20ABE09E870622EBEE3EAB6D30E777F782954125137053E30C3939FCB22AE8CD15C7BC0951B396FB68805E29A8377405170453FC3DC7566C66577;
localparam G6_2 = 2048'h0ACB821C851F8674E22CBB114B84463F4DC0BDF6ED61AE530DB70AC16AB8A34145C45E92421E2476C48AA5346380521685FEBF9280CC256EBAF2185B5BAAC8AA3EE763F3D1DF73E12D839B591C9470033559CCD11D99071E1725BBDF4F3DDD876CA09E63D70B78242577834A85C7EE6C28AB5CFDC87BB8E18D460BB4A489312D429078A8C8757C7983E306934FA7E7F300AE32451B42E6052C5EFBA409F87DEA4307DA3A1CD1443A333DDB58A4D9A60CD488994D421F4A5124A6B4E46E31728FC72BC0004C4A198847195171044C5A5BD3886454C3D2AF1555A40A9E9E0DB79936A808874F3C274EC6D97C75AC31A90126B901B0062F6B28E8B9A15646228783;
localparam G6_3 = 2048'h26664A6564724DCB72414202E6DCF1E0050134E43544C2BE1F8E5322EBA77DFAAEFE9197D30EA645131AC9B5A4E95E095C7C82E3FC99B303DA862606A8DACACF4253046B856FBEDC9FE8E54A03A2706445BB99AC87EF3AE340A0A87FA0BC0825125A82FA498CC5F4BA011AFD11B7FE689408479D931C75F090615EA47611CB3A60DF87AFEFA745B4D7196A0ECF1FB4C996FCD21F9690C178F99E2C6EB78F8F5C24107C97B75FAE4884490D75C1948F24011729D94E335AB63CD6BF5C072B7CE9DF4C746D2A9665F4CE35C35EF3E82687A90BA2A0F1172B35AD55E16E5A572340B92463BDE5A646C9AC6913B3477D6A41E1F1DD27DA6A4D68B9F605510ACF4DDA;
localparam G6_4 = 2048'h1008CCDFDE977F1BEEAADEBB60840DE368EAEF98F8F989CE1B4726716369366E9513B7CE47080E80CA553DF348C9CA0DA777211A6D8796347E4A3EBC99F8CB00FAC1CC3638D75AAC5EE5D0A5C7A7B14DF5AA51D545470E8FD2375379E53B974DECE9A74A8968AA6670013EC96AAB3499A9A5DED3B628AFAE56C6A56091854E235C085E03B2602C717F674F68DCB97FE72A93FE745A0C7C9869729CD88C3E6F6BB72D10F07E5CE28AC636D01A0123C82AF30EFAB57D08442BF4EF07A4C6D27F0D14B13854404BCEC54E936C6365C42D5E9DC5614BE3F499577CF743EAFD02D6BF6AC0AF81371696D2F7A72CEBCD5808A65BDC95BEAB90EB2F56EFDCB3AD63C008;
localparam G6_5 = 2048'hD5A7748FDE74A9C1520A6A4953763CD925A4F13D60E9E6AA7419900A9B25738D68F6654527B4FF506BB862F94E655FB7DBC7DFE25757D89E64A04A183BAEA52842C5664B2BD5A8513D34ECAE5A07B541ED53157FFC2EEE2D4904ED512B7D3F79E7E61E1F9188E45469C3D164057B5E1EDC7C22147C230669D25CEFF05EF267CC4FE2214E1636CB1FA5A9FD15377088D9209CF4487C52F85A239887FE755AF8CBCD1C1255AD7E4F4DF22BB234503911AC560E5342B8C2D8E449C0D119012D9FA8FEA89F13F92474C3057ACC8F3F2F37BC222ABC6DD2C3AC32EC64C9E28F2BCEE18D8BF8C8E7022BA2E72F4563972BA74A386063A35B68EF730431B2F50CD09D62;
localparam G6_6 = 2048'hA209F1E1AC6A5B6E84BDBFB3D03F4D4EF92DDE9266804A7FB7C2E1BCFC1FAB59731FDD1D38BB454881357E7E3393C7A5389B0CFF8E4242830B2758528DFD5EAA9043BBBB2F23B951EB8C38A7A6D46B5373C0DC9364BAA792EFAD508EF44F9A473237FD9C3FC1719207D8394AA7F039526DFABFD2D066B4423F5E04D1F4536D96AA70843D0E644A8BD5B3833AC64B008FB8159B647279A8178F32CE78E0364DDCC97EC6B8A4012E97F68607F94C62E1878ADDB6FA3A14504C20A434B3D01006C860BAD0993BA9C39FF757F139D9C593D921CDC027A488B41DEBD2B3A048D4BF88CDCBB7E42DC6ACF9F01BA066837263CAEE3E24BE80563A2072D73070DD93CC22;
localparam G6_7 = 2048'hE89C9D6CFED0EDC9449329D2E825A419F75A9E59690C5A49AF243D79875EE3C29DDD237342DBED98D56C459D1933356F7C7E55AAA551F52DC042CDDBA704230B4152D16265C111E43EBEC17637D7494C75E9406513706FE4E6E6EABC6B9A15659D3D96D8C0580697F3A62A8A492DCFE7EA558226C774270EF3EF6F4613C3A9D07A5913F602BE94ACCF670FEE5D0BF728BF1B98AF8D1416838DDC7DAA1D5858D4B4E0E642275230DC49E15B3176309AAA8D61B519939287604E2FBCE2E4A2F2AB1794B9CA626B519D69EBA4560D10F9D707E08A3455D272E2B308E2A41E2879F528B32B11BB5B020F2421427639D1B47BA812532529F70193E6E12A943257765F;
localparam G6_8 = 2048'h2999ABEA7B201F23D23177B87205706E8BB213E4A119A1A693BC3A9418C207BA3038014F4FDCC1E16EB1B6B51CDB57E22A94413D822E43CF862EFF9A6AE4E46DC3142548F1507EFA1381CF20CD12E77C42C2456FF57FD6DC477EF74B6A95CD971EDC80302E243E4EA9B243A469ED782634A8A00FCF9F834CA58CE5DCFAAB35574E8358D19FF1DAC0D241E96D3F3D2565C34B2B61521554CB438052A28D97C69F3D14600B240F7F32BD98E93C190AF482E8ACDB4FC94DA1402370C268EA9B4ADF7072938C0CEA7F799AAB50B2D172C8552244356FC589CBDA0B37AC2D337C3096CDAB8EFA354041CC7395EC025CDE2250D7D28EBB176C16367CC1251980F30DE7;
localparam G7_1 = 2048'h1BDD4D3BF61638FC3A34176129C3365B89984BB503EB2D9CCDD267D80DA46BB81446B03B1D3EA5634AD28425FC1C01F19261F3E036FE803B705E2AE708750A8299DC181652F2D96AF20DE529569C1BE6CF428ECCB60FB5BC8D1DBEA898717EBC806617CF9993A6CC867CEE9DFC5F842742E21937DC2C41990656CFEBA5C2B242C467B13221B3FF4C6FDB8D0E0C531E5B908D0FFAB704286A1B18FCDDA9E4DB68050879A95CB98AA830346B7C5B52EED792294B4A454D93AC0D9D5651DC20CD25165A582027861AFB2E5184D60939C546F88B5E45A45ADC709D6AD83C1BC613E6DCA133921474C6EF467C15985F95433CBA23F0A70185E8331786FCB1E0B266F6;
localparam G7_2 = 2048'hAD91F64689A3D5EED9B082F14E82ABBA79B6F153B4D8180D405ED02D10F1F7C21C6D3A3E90F38C6659118BE59288A22D70566799C9DA6DCEE405375F1687B1BAD508490844803FF71F895F9CA6B980C45D650E73DC65D5F08A7248B8E25C2EC8C51C760A61BF3141F5E593CFE56CA78187BF222DB8E923E404E1637C75B75232486C5CC517E2AECD324A673AF4C460A7C91652F953D5770DF4073C3E488A21DA79DDDA3209C146E2B877B7E3442BD7CFBCF762AF237D8DFA35BF900D16C30A8A87E5F8708C2DD806C3AA75219CEC757AF42DF8EC1232B92FC304EAFC94DA86031989F013CD040CF6EF8C81683AF6CFD8595C424F96FDDB276E61780197EECA4E;
localparam G7_3 = 2048'h1EEFD03EDA4FDDAEB2BAA42219CCD8A0EF177B4D18B3E4CBE21D7EAEEA5AF3252FD3319915BC6D01DE37595EA78A16D51A291CD2FD3FFFA2E5A34E71CAD01AA5287A47021ED6E2AD6621656CAF530476641E150DFBC873EBEAF56D335DFB1EBCBC8EF0C033D6E1E020C5B49839390B2EFB91BFCE7B9388520DF8EA6B5151812B593D9BB0A78927408C2CBD4986ED59DC8793C4D98C6F70657B8B86F4F29DF6EC20577C05670398A9152CDA2DB99421D39E437295DAD244203200A93FF3704DDC87CCA064E43FB6CBFC93FA1A795D225E5B606E8CE719EA9CA4B1B35F51891077394C0EACFF18AF61DC7CDF5DB10BB74E12723E2C0BCA0DFC8F521769EDF068F5;
localparam G7_4 = 2048'h76F11C5C1AB8B5E38B41CCB819AB5AD324C786971F4AE4DB55FF8BBB60216804D3DA940301096A9EBA152D5EF838BE3D1C31A72391D7083AB89E0E8FFB1F3E83917D39F9913464C6FA21E781CE5176DEFE7187B9A6793BBB8329EBD27BCA1F850A45974B9D0074E8A704D866BF01A033C89E49A7AB88C439348FC2610040B59A4FCC489AB3E9C0713CF39B997DEFDDA8CC5D03F1E53EB2EF8463B9BB9DDD3CA3D13A579AB1DA3749E4C3A75B553992053FE9BAF9B1B9524F24E7BF1992F50AE8382A8E83D255B7E1B8FF4499C79A4633B09806D36232FBECDF7D7E246265D9E4079E158D50A5D3B163775EB3E9ADE4CF2C6C7079751BB46D70D38DCA193C64F0;
localparam G7_5 = 2048'h0B9712BB220996574F167F9A7AE52563CAD84015909668AC1F55C4C0719779D55A80BA0A542836B87E510B450DBBDF1E21A8212AA990C3575A9FA0AA1A178F3DED7B2B10C597D33094091BD7565C4052255939C63A9FED055B8B0AA5887A4B8E9ED04FBC17EB17828EBC46D5A934368D4E031A4BCB704814B5E4E8C2D9686D438E8B9D4526E172A5B1A88C319EDFA521933FD6E946477BBA0B28DDBC1DBADCBA94F992DAA56C0902709109E26678150F7E3B5E2E4AA0B14A24B80E68E3F33CC01A8C7C7C4EFD58C5CB8073A3A4A5103DE5C758EAD452476E989788733922EB58740D2C196E55C33595796A9F8C57D398DF0AB29E00E5E39EAEBFA95E3A6D64E4;
localparam G7_6 = 2048'h56ECD1DACDEE97BC991448B100B7EDA59741BB45A9EDBB41EA0DE223CD388660F957DF0DFC98843D83D72FE1C29D4E75279D1E2ED489B75E1BC5B2A00F5AA515899506B69C9998D9C1E3D7BB7B84B9E298B7002732D05039D2E93C8435EB7E31E0DDF9B97446B3D97E36DA525203215ECDEF79554CF5E5571CD800F12418337CA7B51AD5374CC84633065F38D149B264A862534D90A46F820519843B8CCC23D98A32575050E95EC8FF76FDEF05DD6A75003A857DF07C55BECBD819B46BD1EE8A6BD5BDD92297C610A2CD7E61205C43A1F079DB78692D244F19443A28E7535FFF6439E340B7F6B67C858A77147AAAE2390C3C92503B7D477EE3DEE36225B19FBF;
localparam G7_7 = 2048'h7C60B988F69CF60980C74B9C3A810A37777A9EC952EC956143ADE443B62FBA6F27271160534792A11CFF0D12C555D17626152720E21A7B33730C0CE49A33DF53FA32091625FA3889A7C302ED446B3CCBF84610EEBE1341F6565C76D5C4F9C509D89CC9A7C2BC08E388817EFC5A12FD71327FD517324CEEF06ADD4007FF05E48F9729C9DE8986A93219EC9C12CA9FAC73A64A1FBDF6B329458CC886299A466ADDE86AE7AD8D36155D13EAB09C87745BA02B2AB3CACEFAD3449713CC8E2833A13477D8A8F2EFB4B0F5E3B46D6E3B3A22548EB6EA870297BF1DD185AD9B7C097EFE94E95CCA96BEB6CDE712B46FDE905B92AD15E63D81A440C388A37E55D0ED1881;
localparam G7_8 = 2048'hF08136FA92E7B6355AA6A279E7C2CBA24992E5D0F1DEABE3F11F99C8E5B5A85AFD35F63886D34EE2CA668F3EE7047218DC38625DCA76AA419785BDA4FBF72EC81461FD9ABEEAE69652B12530A915D397E7E336926812DB675611ADFD47BE3FC1301F2932744D75E7718DAD094FC26AEA3861AE7623FA4728F269E06BEC3714248616A4B41115E845E4811D7B6A35A3414EEFDA03E21E522A71D768458A4D9B7BF45F01DCCCD53F5FD5FE95080DB7212F58E9B1E7CE060865638AE7B71777D90F9CD45A6B0082203D308A576554861FDB46BAB3D80B31397A5DFE8673DEDF435433EC3A455E6CA7F7FC7E6E24A731FCAF458C81F38626915F34A41D24B338CAA4;
localparam G8_1 = 2048'hB2B8CEF1A9D33009BC6B916CA440C7A4DA3EC4BA860A497168B40F8A2762012EF52C3554F3C1C5B14F8CFE1EE22EAB9FF6447E1D86FCDFB61B40B9CFCA6A825929FCC7C74E63B107D27A9749E21C8C9A8D443CFE39D829B5000E17871A38AB90199F76EC9BE0A377782C5D03E14F9D1A548BEED0F963BD4B61E5296AAB741D699914496B4C88D22863DCC7C8C225624567D36526D30306EE756207D9F8750DADD642EB8EBCEB8E74270CB1A86F8EB8D1FB6799D04C5B7F634212D61762ACB95FE77EBACDB131C84664503D134D1F13BB1EA5D8DFF6BA3A703C9E91D46B532C8FAB2F9A547BF24BB1DCCBD1280AFA889310B9ECE9B92FDF8FBA1ADDE0B61EDBC0;
localparam G8_2 = 2048'h9CBACDA8BD56763375A13C9CFE14E749DED9762784D968464354A7B8E635A496F25F3D6E298E7E950CDEEFA2C5919A65819D2FEB946179E24490621955EEC9822CB8698BBBDDB575969A734EBCD2673E839A2D8EE6CC8FDA6A55A05DB6FA9E68FC57F8F854348B440F47C8066E5A174301B934833DDBF0F4B989FE6C4B33BDB2B342F3E5A0355BC96B0D0718DB22FD1309E0640F2287B7BB152345C5F07AADAF51FA0127CF70BBA3CC1E78C3F7B41A069A0E8DC8E63348DE0A593C25C2546A85427EA20C48DE36E6F04256E181CBC0E269682DC525980D47E8B38926ED527E6F54B40A1E923AB9CEE23935C7EAA99071C27CC7A6EF14E177A816482705531735;
localparam G8_3 = 2048'h5F791CD29EB3892A43AC636F1F371703FAFD495D359CCD66165DD93D40B51E9E5C1B118A2AB56BBB67B0BB0BD2BE5A6E0E636D5C2EB8C32C312739E1C198F32E0C9DB604F717A2DA1B41684961CD847C005FAC40623F8F2AC73D6CED71F89FC8DFBBB8E10E571A61889685E85632308CAB3666A1EE07476647D1FB0ABDC4F43744C5F07B5683463213B68366D49EAD2B55D02496806F50C8D741142130D412D3727E94F190371284A9D8BAE431E01CBDD2BDA3192C9B4C90A96444A555E3BE1DC0CD5FD5BEA4EC72BEF93990E9D256104E2C124FA9C4D9324C85DF12B9FD0F9401AA477251184E83E840DFF30347E511D07A13083F354657A7BED93DCF3965D5;
localparam G8_4 = 2048'h9C25BD30B35F6EC38FCA2AAE1B45AA675AAAF4C1298F679A44F550DA627FCEE84D0CFEA9CA03BDB5919AAA0F3FBC5D2A564088C14AC633FCEC470CF0598DF1ECC13B042617EB5E720E368F39600E5F0BB7B6E9B3F576C223945B0729B6BB212771FEB035941C8C53C3C9CA3CD2E047BCE2382CFB8EF2FCACFD65CFCEB616753FA507B89CCEFFE8655B1C68838D6DB571B3C909B51CCAD4DE41E6040025970E672606C28BEBF7C55E95CE9168AD3885DCF0FFBF2ABAEE45AB93ED00FFD9B91F2EF6B235652ECE6B93A7F5B538837E7EC0F1570129B2724CF59F9344FEF0AE924914AC9585164A0FED39B993A66459265E3911F83C261E29BCF1361ECA41748848;
localparam G8_5 = 2048'h584771DFB4CB4C32968BD6B7747C7108F6E3383F4BDEEB3BEDA7F7E266F1EE2A027A291AC4725AD3E3290A7A4567B018E983CEE155ABCD9A6F2D1489AFD01E3912F978775869CFDA5F029BAEFACCD36D0C7670C767156E15A767A98A96F4FDE95E5F84201483BD9870CE43F692C205B5CF1E94B0001A446DF726ED6BADDFE0330E9A0927D8423A754D948AB12F69EC8EB0273D4D4F57366D9A943D59E00125BD9387DE7D332706733B4A221ED46D7CFA0F7AC71FC3FA3F0499A167DEC4E574F16EC07E5C0692F99C4897C835DF3E7658734ED21F93AF188A1554811B47532F0103BE0DC2C49ADD8DF6394CA1C864D7AAE11944BFFCF7351EACBEAA77894F5CAA;
localparam G8_6 = 2048'h8E081968FDD6AE371FCD85FD333CA80C307243464B9EBF24CA01D7F14081DB9C5F4ABD5DB154E0F106F2CC40CD14AA02B33986B97A6736E5D93F10C224BF9928DCCE6C6ACCC7EA37283F12692E5352E86C5545C8B9C8DEBE00B45F9F750C3DAAA92A2D8B65B28F7FA72F08573D3930A46E7A9020128E45B7DC453D6829DC6CEE81C68365166C0B68A6A7FDF67CAA49CA49D4BB3D13D8A4B113190788AA769461F0790560C49D648A5938A3780523688CDE07CDAB3ADAB7F227FC75C619BEAFC2D790C29671481D6888D80B8563B9B29A0CD37F0E99715F2A0B3CF86D05A0031929DC056640FF7D2D4C0C0BD3C2BCEADEE7961FACA479E9A85542D62776CC701F;
localparam G8_7 = 2048'h72B0CB2356D93DD9612B58302AA3838823AB4E6A2C837E5BB153AA3ECA12833C5133970F1E584F7C2DF0FAC943358DF4F04359A2136C0F476F315696526033320194780A7BBD918493F132468322A132C480C7A8D75F28E1BB840C47C0A6BC8B0D5A8FFCABD6F47CBDE16E7873B0DA243AA4EC934D1933232913979226AB9EAE0EADF24A0FE2123F2A907795C778F8DB350C7CF77AFEB04A10847C8A2FD7818600396739AF95F87116519D9F2A45718C8A6932141C5E6F0A17F4FB381E32813C1418E424DC60C9BA1780B4726BD67E3B71A13B6631A6E0C268F21431A9CC69B17B118AA6400EADEDB49BF9E44EA7FCF3A009AF7A88323866EDBA6CE6A7DC0807;
localparam G8_8 = 2048'h93B6B0D8BC58456ADE6654F69510DA2E566B8AEB86D6AB0C3EF02A4D2231B446CF8A04B0CCD0166C34D332F0BE496504390F439ED900E3D45A77A6BBA9EE9F8B7D61A9D65BB7AFF8EBF71AD16F0C2030485B86BA296EE297085D7E231EA5883EA227F6013B89A6E12CBFCFE16E1377A7EE7F9AFBC56721738717D75A25786B78440EC9EA2905E03BBEB97EF70E49552E7F07467FBF40A3031D6DE9ABEB79C9546D5C7D5A927ECB1393764A165EFD559C65C531E26639530FB8781F4B5258DD62EE03F77965EC355324C58A5775F1F7121B4A505FD94371FCF2CCC6FE6689451239DB6CCD16AC89259BBBF42D48F408E4B3DDE6FA3D573EA45E84FEEA1B11296C;
/***********************************************************************************************************/
input clk;                 /*系统时钟*/
input rst_n;               /*低电平异步复位信号*/

input s_axis_tdata;        /*输入数据*/
input s_axis_tvalid;       /*输入数据有效标志,高电平有效*/
output reg s_axis_tready;  /*向上游模块发送读请求或读确认信号,高电平有效*/

output reg m_axis_tdata;   /*输出数据*/
output reg m_axis_tvalid;  /*输出数据有效标志,高电平有效*/
output reg m_axis_tlast;   /*码块结束标志位，每完成一个LDPC码块的输出拉高一次*/
input m_axis_tready;       /*下游模块传来的读请求或读确认信号,高电平有效*/



/************************************************进行LDPC编码************************************************/
localparam STATE_waiting_data_in=3'b100;  /*等待输入*/
localparam STATE_data_out=3'b010;         /*输出信息位*/
localparam STATE_check_out=3'b001;        /*输出校验位*/

reg [2:0] state;               /*状态机*/
reg [$clog2(n):0] in_out_cnt;  /*输入/输出计数器*/
reg [n-k-1:0] g;               /*生成矩阵当前所在行*/
reg [n-k-1:0] check;           /*校验位*/

always@(posedge clk or negedge rst_n)
begin
  if(!rst_n)
    begin
      in_out_cnt<=0;
      g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
      check<=0;
      s_axis_tready<=0;
      m_axis_tdata<=0;
      m_axis_tvalid<=0;
      m_axis_tlast<=0;
      state<=STATE_waiting_data_in;
    end
  else
    begin
      case(state)
        STATE_waiting_data_in : begin
                                  in_out_cnt<=in_out_cnt;
                                  g<=g;
                                  check<=check;
                                  m_axis_tlast<=0;
                                  if(s_axis_tready&&s_axis_tvalid)
                                    begin
                                      s_axis_tready<=0;
                                      m_axis_tdata<=s_axis_tdata;
                                      m_axis_tvalid<=1;
                                      state<=STATE_data_out;
                                    end
                                  else
                                    begin
                                      s_axis_tready<=1;
                                      m_axis_tdata<=m_axis_tdata;
                                      m_axis_tvalid<=m_axis_tvalid;
                                      state<=state;
                                    end
                                end

        STATE_data_out : begin
                           m_axis_tdata<=m_axis_tdata;
                           m_axis_tlast<=0;
                           if(m_axis_tready&&m_axis_tvalid)
                             begin
                               m_axis_tvalid<=0;
                               check<=check^(m_axis_tdata?g:0);
                               if(in_out_cnt==k-1)
                                 begin
                                   in_out_cnt<=0;
                                   s_axis_tready<=0;
                                   state<=STATE_check_out;
                                 end
                               else
                                 begin
                                   in_out_cnt<=in_out_cnt+1;
                                   s_axis_tready<=1;
                                   state<=STATE_waiting_data_in;                     
                                 end
                               case(in_out_cnt)
                                 sub_size*1-1 : g<={G2_1,G2_2,G2_3,G2_4,G2_5,G2_6,G2_7,G2_8};
                                 sub_size*2-1 : g<={G3_1,G3_2,G3_3,G3_4,G3_5,G3_6,G3_7,G3_8};
                                 sub_size*3-1 : g<={G4_1,G4_2,G4_3,G4_4,G4_5,G4_6,G4_7,G4_8};
                                 sub_size*4-1 : g<={G5_1,G5_2,G5_3,G5_4,G5_5,G5_6,G5_7,G5_8};
                                 sub_size*5-1 : g<={G6_1,G6_2,G6_3,G6_4,G6_5,G6_6,G6_7,G6_8};
                                 sub_size*6-1 : g<={G7_1,G7_2,G7_3,G7_4,G7_5,G7_6,G7_7,G7_8};
                                 sub_size*7-1 : g<={G8_1,G8_2,G8_3,G8_4,G8_5,G8_6,G8_7,G8_8};
                                 sub_size*8-1 : g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                                 default : g<={{g[sub_size*7],g[sub_size*8-1:sub_size*7+1]},
                                               {g[sub_size*6],g[sub_size*7-1:sub_size*6+1]},
                                               {g[sub_size*5],g[sub_size*6-1:sub_size*5+1]},
                                               {g[sub_size*4],g[sub_size*5-1:sub_size*4+1]},
                                               {g[sub_size*3],g[sub_size*4-1:sub_size*3+1]},
                                               {g[sub_size*2],g[sub_size*3-1:sub_size*2+1]},
                                               {g[sub_size*1],g[sub_size*2-1:sub_size*1+1]},
                                               {g[sub_size*0],g[sub_size*1-1:sub_size*0+1]}
                                              };
                               endcase
                             end
                           else
                             begin
                               in_out_cnt<=in_out_cnt;
                               g<=g;
                               check<=check;
                               s_axis_tready<=0;
                               m_axis_tvalid<=m_axis_tvalid;
                               state<=state;
                             end
                         end

        STATE_check_out : begin
                            g<=g;
                            if(!m_axis_tvalid)
                              begin
                                in_out_cnt<=in_out_cnt;
                                check<=check;
                                s_axis_tready<=0;
                                m_axis_tdata<=check[n-k-1];
                                m_axis_tvalid<=1;
                                m_axis_tlast<=0;
                                state<=state;
                              end
                            else if(m_axis_tready&&m_axis_tvalid)
                              begin
                                if(in_out_cnt==n-k-1)
                                  begin
                                    in_out_cnt<=0;
                                    check<=0;
                                    s_axis_tready<=1;
                                    m_axis_tdata<=m_axis_tdata;
                                    m_axis_tvalid<=0;
                                    m_axis_tlast<=0;
                                    state<=STATE_waiting_data_in;
                                  end
                                else if(in_out_cnt==n-k-2)
                                  begin
                                    in_out_cnt<=in_out_cnt+1;
                                    check<=check;
                                    s_axis_tready<=0;
                                    m_axis_tdata<=check[n-k-1-in_out_cnt-1];
                                    m_axis_tvalid<=1;
                                    m_axis_tlast<=1;
                                    state<=state;
                                  end
                                else
                                  begin
                                    in_out_cnt<=in_out_cnt+1;
                                    check<=check;
                                    s_axis_tready<=0;
                                    m_axis_tdata<=check[n-k-1-in_out_cnt-1];
                                    m_axis_tvalid<=1;
                                    m_axis_tlast<=0;
                                    state<=state;
                                  end
                              end
                            else
                              begin
                                in_out_cnt<=in_out_cnt;
                                check<=check;
                                s_axis_tready<=0;
                                m_axis_tdata<=m_axis_tdata;
                                m_axis_tvalid<=m_axis_tvalid;
                                m_axis_tlast<=m_axis_tlast;
                                state<=state;
                              end
                          end
                          
        default : begin
                    in_out_cnt<=0;
                    g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                    check<=0;
                    s_axis_tready<=0;
                    m_axis_tdata<=0;
                    m_axis_tvalid<=0;
                    m_axis_tlast<=0;
                    state<=STATE_waiting_data_in;            
                  end
      endcase
    end
end
/***********************************************************************************************************/

endmodule