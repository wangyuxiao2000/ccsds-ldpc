/*************************************************************/
//function: CCSDS-(20480,16384)LDPC编码器
//Author  : WangYuxiao
//Email   : wyxee2000@163.com
//Data    : 2024.1.24
//Version : V 1.0
/*************************************************************/
`timescale 1 ns / 1 ps

module encoder_20480_16384 (clk,rst_n,s_axis_tdata,s_axis_tvalid,s_axis_tready,m_axis_tdata,m_axis_tvalid,m_axis_tlast,m_axis_tready);
/************************************************生成矩阵设置************************************************/
parameter width = 8; /*支持1、2、4、8、16、32、64*/
localparam n = 20480;
localparam k = 16384;
localparam sub_size = 512;
localparam G1_1 = 512'hB3538BB9F7D8270F6BE80736B2F204D0C63A9A2024357CBDE3E390021DA5C95962AC8FB8A369B0E17A4714E6210F9D7D0662BDE44BC3779D2C88BEF3E44813A0;
localparam G1_2 = 512'hB997D9EF6DD0EBABB63CF71B9EE59FE8802CB1488CEFAAB78E3510C7FEDAA8C398B27F71B80AF19DE9B0381E53941FAFFB4707D29BE7FD52FF8F6EF442FA6B67;
localparam G1_3 = 512'h9A71DB5B2889C799A2BD40E14236F3673F0DB3B19BF3E300B4E383C0C16BA83803C0D716DA96D9403D5C1C49BEEACF710E112CDDAB515D434F639F7B0633F35E;
localparam G1_4 = 512'h25EA0A723D9A66F247E31047876297E68E27AD4D50F814C974B7F268C9AB9CAE6830C7DBFFCBFF2FFCAF7A530FACFC29ED8EC1181AC767344EF7FED03A18AFBA;
localparam G1_5 = 512'hA6F5BF1B46D774D61759C0156846CA20FCBEA4F233C66CC2CC50925A9D382ED80CE05657BAAAD936F33EF5DDD0DA7E194A5E61171C52EFAF0A709EC7DE180B2A;
localparam G1_6 = 512'h3577D80F55CD833D6335A60685D48F7612385FC95934AD61E2186AD3A4A9E97B2B76E0FAE4047B3E8819B1D329CA462DCCDBEE2C6462AB140563FB2AB5268752;
localparam G1_7 = 512'h12091D2DB3E059342F2AC97A72EDA24076AFBFEA745AC6B833DF6A79ED43BE1FC0EE1DF1A137E31F483087C797F46EA589E2A5B5683636102B9C3F28194197B7;
localparam G1_8 = 512'h972CA2AD1B9AA59DD81548046FB0717C89D7EF650737B8A08864F02F895217617759FDC4798251823730518958B57B59BE1759CB3E756F3BAB41EF2FFA4A707B;
localparam G2_1 = 512'h1E00934830FCEBA8C62C00CFFD779FC2004E253733DDA08BFFF326AEDBD7E03FD4B4032B0F2B364FE9E9ADABD266B9BF86551E0D3D2515AAB47E660C44E96438;
localparam G2_2 = 512'hBD838E264AEDABEAE7500274CFEB5E8F60B908266198DBC8FC93FA1FFC7DEE2942FD59A3F7C732EB9658FE9C64F1BED6A0F73FDFC04ECE9B70DAC0B988122C8E;
localparam G2_3 = 512'hB00D259CDB47FD148322C347368DE8620ADF687815BCD6CBDBB68114B4064ADAA1C857644FBD5894D48E2EDA5C977E46CCEC7B070362D9DA3E1976033E44E40D;
localparam G2_4 = 512'hC198B44DCE89718691F9E75D505ED4DC519CE946C0C7BD6F0158BEAADD055A4A4FC4487B0CA393FCA3C06DD1A80F8C76FC033922A6261E62F37B0B323EC289D6;
localparam G2_5 = 512'h2C157C4FFC4FE9758491D28C767223F26969E440B6154B2BAE49E99823E2358272B8E83451BC8707D9A97B88B52537CA00CE6304BC85AE88889AEF1058D9A576;
localparam G2_6 = 512'hF7EF1D9B1286D5DC668AB7FCE17B7FA055DA8517AE35DF8AA22B183681B1EA070B3A909824BBCE4F0EB1EE0A7DD64AF8E6C6B066816B2C575784B9C7354FFCCE;
localparam G2_7 = 512'h4E1BF3AA8165566940AE8A58D56333A03C35187597BBFE2FD8961DE59E362EE63B3F47A92545CC797C7DC1A2EA2240ED45A2BCFA817A25EC1375F745DD8B8F5C;
localparam G2_8 = 512'hFC92C0B6E992E2AFA1E6F0D726262AF42DCE9707D384D5651566EC07E92EABF0EA78B71A22CE7A03E5A1FEB0EA5B9091210AD96B898E45B4B8BC45B6468CB17E;
localparam G3_1 = 512'hEA8C74DD4B365B5EB3A04D4628DD782CD7F46BD378638D39BE6216458D35892847AE2DA6F71D4B9A7B1A7AF91EEFA9674978672D401B7C208012B2649127C837;
localparam G3_2 = 512'h07C5C4127373151592FACBEC45965DE9D17A0AFF71E32F844252711A68EA359EF7E30C2551AE8CE8D1D1D6E9D8F4D153D0EAA3A81AB252F44AEAFA8095AB56CE;
localparam G3_3 = 512'hA043F3010FCA8617EC9EE4128D76AA7DC0F949D5D48DA530E71973873064E49834EC4C661DBD6D50F2E54A55E0155F9C2A4B1C4A9DB61283114DDF6DD66BEB39;
localparam G3_4 = 512'h2F8253A507C913AC7D91436A5388372EA05E6ADEFF988E064CD0FB1A6C3C96F128911DD157A93A3038D700272DD7CDD62ABBC98D4E98CFD01659449315BC3FC1;
localparam G3_5 = 512'h976D878BFC6CBD2752CD8C77D36C236457AA7906F6B9AEF7704130342786557BEEE6F8967FEDE8C2ABA74D1576E4107EFBDEF30A22439B338EE55BDC32F7AF10;
localparam G3_6 = 512'hD9D124ED292320D29419EBF83F29D619821B6D798281B8D216BAA908D74C29BA3FADFD8FEF430221A81572F4DB7BC78CF73767D44D1C1D334630405795380A76;
localparam G3_7 = 512'h360E71CB6FFF406AC5A4D60C74F4490DB721617919C640DC533EEE2B05D5D13ADD823C1F2B00FC4512E661EC73B686FBE73A9EE211B5FBC94C311648C539C8EC;
localparam G3_8 = 512'h0116286ADCBFA039876252D53449E1155F754CE4813BB2DDA3A76BAF503228909E989EDFB66DD52CF9B9AF7105F49360A9BFECB3C847A60C9F826237C66B430A;
localparam G4_1 = 512'hD06FD1661A0D12C5438F5B7CB27CE6CBF1363F23DCFB9FD5A260F1B71EBAABD770B48C3D8F2B5503923371D2A09E028EE17179554599A62981932E0FB6A9546A;
localparam G4_2 = 512'h68DD5428C5D0DE1710A817EE122FE2CE0B436C71D78FBC069A0080B0EFFB9C5BB9B59D46C5819BF505D4370AC83AE69626A2940C6609280EB931B50C4CD34628;
localparam G4_3 = 512'h3E0F0AA4403BA786C0274681EC0B120204D123A490422DCA34CD2CD8FB205039CA473B624535148723ABB72D052100B3AC860151E16EA11BCD6AF40748B2DF32;
localparam G4_4 = 512'hDC18EF57734121B1882DA0EEB9AF79CA4960174BCE22F1F4A2C48C9C361ED85E1AE78B16A52496E31DE2C2AB6577B9093A03749A02CCB80D2E5D81624723C9DE;
localparam G4_5 = 512'h3351927BA5ED5F34369A62E64FC5EA2C9654A21E1D3BF7298950F6535FA5F1EECB28FEB09BDE952A7E91CE5D9450F662E8991B7932C087467BF24D86ED2CBB4F;
localparam G4_6 = 512'h674DC69631CC77F63E115E99B541514725861D1BA6E68F28930B5C7CD806FE81AC4F959D786246CCE8E725E87ECFE8F6BCFF98102284A95B461FF751D6912E6C;
localparam G4_7 = 512'hAC471FE904A7A0CAC20F9159ADA66EB3239C612A2BA314EEE1A65DEE50DFF1556CF5CFC4B1B7210F99D70AA7A7C8166D0D76CD1AC2088104AF87658CEEA573C5;
localparam G4_8 = 512'hF1BDD31317E7D65CC6413D2E1FC01F2357F1183377545D455EE12DE65E9F51AAE7D01D5315AD8A02B54416232B18523765A70963BD9D0006D08CEBE1219FCC0D;
localparam G5_1 = 512'h8420292DEB608258513FB910A2F0F49CF61197ABD066F7A0AE210E32ADE24262226E6BD13A1CEE00C5794444E9E2504412D7618C63BD5534E7042ABB29042963;
localparam G5_2 = 512'h16C511866AC1EFDF8FBCCB01BD9398B23144076D85FD79FB68BC9BD61699B867CBFD5FE5C2E6E835ED0CEF0A59891CCE0BCF18CCBF7C0F7886F298E46B3A8D07;
localparam G5_3 = 512'hF1BE8F2486A7CA53A54EE787F890E9B505A5968B5A6D03223F8759768972DF1A0D65178CCF8A8F4D0337829C2432B11F669046061CDCC347B30E5868D7B24387;
localparam G5_4 = 512'h6E019E4B229FD71B69FC313374B42D6B44BAE71AF738499C6BE8ECD5D709BB57928C5EE4C318E3A87E031D0AA8197E3A65ADA191B8FBBF5E987B6F550A105A27;
localparam G5_5 = 512'h8C7CF04AC61AD7326F74CA175C7B30648F8784293CA1B1C0D79E6170D3C7A7A0D08977FD393F73FCC4F96E5D85ACAF4992D18D617E1DDF5BE9A73210873BD833;
localparam G5_6 = 512'h86C76BC7FD47A4AA911863B6DD693E9F281ACDD41324253E3ECF9B4E24156ED438E7FCF609910594761BD37BADDAC09EC6A034306DE38BF7AFB8CB1DF5F7333A;
localparam G5_7 = 512'h1E8D1E73CD7B81A0513875DD7DC0F3A589CBA83E507C559E444E6505D200F05B878EEAC789D44690CB83289F0BC4B11F404A5A812A6DFE5C252BC4100CE744DA;
localparam G5_8 = 512'hD2CE4F2EE99D55F986659304784B6C4F6DFF8F5122442355A2934A54BD4DB552EEA5E144DD567E45300A268C572ACA4EB01C71F246C1F0968BD66B2A71A95550;
localparam G6_1 = 512'h975CED50A31C625C28A5DCB0806EA8B42655F38F9F3CC859D83F0DB9670A51B20C3DBCAF1BD42C03D303B43FA30534AEAB5FB9A591B34E6C758D881429F63BD9;
localparam G6_2 = 512'h1E2FA684E31F67C3C0D57210639D8CF97F245B17F9C17AC4A9A456BB21A20647F1CF4BECD10EACE7CE3BF0E6ACA14DD9A593593BBC1FF465DEF93E34F20E14B6;
localparam G6_3 = 512'h55C932C07442525E83F286AE86294812116ECBBC7CF57AE60E182E708FD2D9FCC58D38FDAB79A3605935B1888711E4674BA85EB3E29580A49EC8ABD194755ACA;
localparam G6_4 = 512'h94475FF296EE5C7C9B59DF29C6E890CA74166FCCE2A80E7F43670131643949A2767B9F8140662259F1DF87721B22B93F188A6496AFC4259B5258EACB459880A8;
localparam G6_5 = 512'hBE4D2F12ED5E1BC2D31101FBB6DCAF257669AD2AFC871DEC90390C9F116E3AC4538F5D55771FF55EBC6C2F4802602A05A0B00E5703FE062D712B286BCD776B91;
localparam G6_6 = 512'h90DCE859CA64B5BD916E4218C52FCED93891A379B27C45195F36CB4E8E395601701E22772316B4F5D688DBD175826F37D1D1961A22B055510F35FA5EF7CB6651;
localparam G6_7 = 512'hCDB0CE2C7C6FFACAA9BEF3979BA080FE3F85DACE07BE3AC8E74DCEC56BF4A27C4E20BC64C3657129AFD1578C4F337F21859ED1F60FD5766564FCCC5047105B82;
localparam G6_8 = 512'h5803B496A6440897359C7F581E34533A1F64898A88FB15CCB253DCAE09E6EB02F72C0B13D7FB0EDF78C150A5EFE100E7045DAF90C0AFEEA4A6DD7FC38A6CA5DB;
localparam G7_1 = 512'h134C3A7C95EA7C5AD442250506BBAAB9D1A601FDBF3E04F08BE67958667DBEBD06DB7D7A02035DE81973FBCD8ADE155B9B9089DA13E31E1EA1A97670EFB11243;
localparam G7_2 = 512'h2F404C0EED4EC9314FCFA4352825E6A168861F06C72C245460CEC14D464FFA5EB780592CEE2A2BA71D0C67E88DB57B5BA3DFAE45931E51FED70B3BA3E4B6649A;
localparam G7_3 = 512'hCE468279ED2FE97C99EE078C09FE40655A0A17910E87550AE7345A2E9CED29A67AE31A15C586079CCEB46A907393BFBA1A7ED80641C2C5A2ADEC39994CC29920;
localparam G7_4 = 512'h8F417B71196A084C18D8482CB1350C709B2A5CB6411753330755DE3E6E90D7613BF7D9AEAA177DA7E3C1E55D7F9FC1AD86BEE86B839DD7B7129A37FEA0B6B800;
localparam G7_5 = 512'h888A4F502A955E927D97929F50C17773C8EC54DC1113832B153F1AB7AABDC79B0C07BB03F65705A7DD79A20711EF9B5678749A609106784CD8F65010B0B79CCE;
localparam G7_6 = 512'h5DEF02DDC1F3EBD923B45C0D62681CC54E2B353ACB7AFA2BB0D2BB9F6955D54F35AC891BAAB73E9FC4799B0F9B37F7D134441D717884CA42D03DA55AD06CFCDD;
localparam G7_7 = 512'hC93D849E9BAB3EF47B72A29E27EBC8C1857DEA14D78557DDFA8B671DF22D38A7B7F22EA14263C8FBE346FF23BBA9DBDE7464F31E6970B52727DEF3C079FDF8DE;
localparam G7_8 = 512'h04A3AAE8ED52C0D10951447AAA873A46BBC80FDF9B1FD6AA51520EB3A7B3FAB8A54A4EFF76A635189829F3757E9C1DD1C4DE154F52B23E7F9A18B6E1CEAD9AF6;
localparam G8_1 = 512'hFACA9EE556665B287EB6E2F50F3C8866321D57F1F3E91049550A0EE541EF5533ABED5EAB92DF594865BEBF5EE39D112AC10AE42CAFFC4215D3802B1D9F95EAE0;
localparam G8_2 = 512'hB21C29C36CBA4F09CFCD9856031FBDFDA4B349B277ABFBA8277F5ADA81D2A2ADDB66007BF92B4C57ADCACBE19385A35ABE0FD30B2C8A8B504F19794C4A393C3E;
localparam G8_3 = 512'h228D137596EBA4ABF53F7A7C5FB07B2B36B5A5680E2EBDBD86D866B4E2CAC41E88FA9A822727AA1BD5EE98E14787929E6B0C5D04B5CDA4F1DE99276D02D25018;
localparam G8_4 = 512'hF65AD93A31924422812734C0B472D3CC0134504C98D04BA4B43E253A084EACB61C9355108779C42A47D8550F95B4CEBF3336C311A5CE3A79E4A6CF1B36458BA2;
localparam G8_5 = 512'hD61C0FD3657ABFFCA8A3638DCBC8F790543FAA5668FAA0976A2D790AB44F2F68EA36A420406A5A38BFB3677BB6468BD01911C389E33137BB264C0E1E4E513E6D;
localparam G8_6 = 512'hFF3C369E6A0CEC9585619045E29E1E1F662C456ACE860A9FB224711802D3F27A5B57F5F8EE59126AC4B5B14C145D9F10E152BF4CF2F5FEBB4B7FC3D255BA0D19;
localparam G8_7 = 512'h961BB2BDD709FC33E8287CAA3EB533F752DF958A891A4AC88242363195FA232D3A224C0C4851D3A0A9C1C5CE3B313DAF8F4EEDE2C5721202A62BB8081639D73F;
localparam G8_8 = 512'h4383A87F666093EBA10DF226C63F0A581F221DF5CBF47A1AA733692ADCE9EA7A02C34771E30CD0266B7B9893B633C2D5964133428AF1EC4172E195592475A82A;
localparam G9_1 = 512'h57CDBBEC6A263D93FB3BF67B5BD5EFA8ECF59CF2FE11FF60BB496E6A5CC13ABE7DC4377A4B86437386CF6A5584AF1DC433BAF671B658662E5B99A8D7286D9B45;
localparam G9_2 = 512'hBF9D7C32FD40E2D3BE6B24A49D04EC07C61450B6CAAD0CDD413962BA16EF75B7EA309CAA7C627218FC3166E4A37F3A3B672B257968A6C6F5E381B2601D47B604;
localparam G9_3 = 512'h5B7C4F0E77E3838D54EDC5087EBC8E89188AB658B05AAEF271E6971717A0C433C6574E81ED3717666A7ACAD775E1A13B507711CBBE50FA8262FE1A009A31685E;
localparam G9_4 = 512'h5C142B773C9FBBA213C48496C4117C0A2EE38A2B4B69DDDAF130D818B55A4B9278F3860BD66DB40D59282152D8746C71B1CA0CE9BA953559387AB3E7205F3D33;
localparam G9_5 = 512'h8D427F23224A29FE054E163F210AA47213884347ACAFCDF9BEFCE88443CDBEAE8158BD41D9DE77D56412C9593A424B6269A73CEBD348D98F759E8DFC66614518;
localparam G9_6 = 512'hD8914D06D54A7BC218D48E785ED4FDAC1E81F9361F00D8DD60DA74ECAE5CF739D4CF487FE04895C913FDEA84B7B490474BBD50B4A568FE75FB1FF78EA6183A9C;
localparam G9_7 = 512'h6935AA7F593F3B99271823E96D33DF922C55711C4C9F149509235B292E3158C3E462DDD674040DFDB36708F0F7CCAF835FC6614600EC0C78F2246406BB01E3F0;
localparam G9_8 = 512'h7C8257670A2A79DE3DD997BFF6AFF58DE9FC0ED0FC474DC357EFD9D270BEA48739F3B0BAF71D4BE6372BB4F2DFD5F25EA59BCB03668C587EC944391AB6159B7F;
localparam G10_1 = 512'h14EF6962B6A9DCCDD86616478543082E25F0308FD76182D4A166A3E262A7BB36447EB125CFA9B7D985386982EA3D9B9AB6BCD1D330B232ECD397129C392FA3BE;
localparam G10_2 = 512'h261E252C76EF048D69627A10B99DA2EC40C8F6574F6991262FDDD271D7F8BB3ED1532875468BC57F41C0A2D77B86684030C36DFD8D5CDAACA2D37B648AEC6710;
localparam G10_3 = 512'h9F11E853BD33A1C5EBB951FCA1D8CCE2DF813BCFE7D10FF701A796E7C5008BA07D7313D7863D8FE2B163A960028A3461D13B77CD4302646BADA8BE843DEDE155;
localparam G10_4 = 512'h3F94F53333D55D56ACB138E9ADFEC1DDFEE0EE286C78790A6E96068181D4439BAED7C42E1A82F6F1889F9F3D8D36EA8481931B5E87248CA0A97E9851DD7A5E93;
localparam G10_5 = 512'hDBB7F58958DE1DAD97A3AD408D56E7A45D902143A6C599D6040433028C977FD1B9071A379FFB29BCB0234EB2E314D88C6269D4D24DDF64C515AD118FE87CF273;
localparam G10_6 = 512'h4616A68D764461BF79161439EA459013FB24BFE53EB822F4D624C0C93ED6DF562B982646C08DB401424EEE70BDE3AE8D53B9F29D1CEADA24D7E6A59E13D0514A;
localparam G10_7 = 512'hFB588EC9E22B6EC02917DD2A656CC48334DC56689CBD2A94C24803D951AACEA3E5B055912F8FD4832E6222C37101EDBF9E74F5D82B34527A79EFBEFD9C33912A;
localparam G10_8 = 512'hC32D7A28F0D9FA4C3F25A4AB87BDC3A1594835BBEE8A8CDA6294B4DFC5C7E67224942079BA4D7483AFE86D0592E562218223EBAF01A671B1BD83F04BF379F7B3;
localparam G11_1 = 512'hA0F38485632B3E3EA87674F47207CEFEA5D18038D4CF5FE2E6118EC36DF92AFB47B946BDEF42750BF1D186F74ECC9AF4E0E94632653FE23E3EEA3F47AAADCF9A;
localparam G11_2 = 512'h5357E6E5C900105FD6F5C1EA0A46FB7F88FE72E4875C03572B76946F7345BA3FEEBD01A4AFC82A586188E6D2CBC78AEAB0D7DE4F1C2B2681A5BEE6E45B66FC77;
localparam G11_3 = 512'h9303F8CA8C4D8CB689A8134DCE8EFF9438312B5B1C762F85F97C23FB1E2D0DA1EFCFE1EA13DE9B8CD254E4EC4949A7DFA3205F0EA1E888AB1A22121F9014CDC0;
localparam G11_4 = 512'h566ABB9BE495337172AF88596F8779887E1501D0276E2A2C68ABAA4D350C2247D4DBE2B29F8B624D75171252C1E97F85DDAF13DE11E7794B2366057982407506;
localparam G11_5 = 512'h431370A6EA73D57F81A3FE9544994970F742D09A5CE768A60AD4058026EFF7EB66B52023989F2EDD3F53361E660EA8B8FF130A148A671F1AD4C65FC8C3AA73CF;
localparam G11_6 = 512'hF15255C0794475B43ED56DEB8138A685AB6AE7705D0D8CA871E94CFCFB22729BFFF9C5A439B7D75B7A9176C08D77CBC2275359BE96F8F47CE3844D1222AD1752;
localparam G11_7 = 512'h6A995821019A29078799039EDB63100136A3B72D784B74F0F888B0D815F42BBDE1EBCA14C8AC9D66690C556206283BCE1EE9065AFE2A8EB2AFD2BEDE20F44292;
localparam G11_8 = 512'hB5FC843EFB0BCAE74536A6298DD0BCF4ECA867814ECF6E67A0A088FD53AB326516FB2375CAD8B9911E53822CD302BFEF8AFD65F83EC4856D7B9056D5A03ED5D8;
localparam G12_1 = 512'h931C21B4945A640824872978623CAF7DCCEA1AEDDCC4AF8CCDD07F38B23C0AACD138BBC4F7CFFD30FDB8225336625DA9026A9EB7545566A246CC2B51A38BF26F;
localparam G12_2 = 512'hD122AFBD41C496813FD598CE87206F0352DB6129EF68F57CDC7BE27A91EA3CBF1BC3CDAF3361632D1B9B81EC10666C1C03DB7ABDA54C36494CBCFCD52AC2FE23;
localparam G12_3 = 512'h36DC5BC3C1246ADBB17E38972F28384127D33A20F846504B3FD3070ABE4080369A953D03ED2A79B19CA2B1DCE2BDDCE0C88CEFA8038000D39ABA55C9391D137D;
localparam G12_4 = 512'h8EC0DD18B606628021D0556D76A1915910C7FDDF1BF1663617C0280F6252F2088AB88F11BDF46F72CCC337C90157EA37071BEFA21AB2A15CEF1D96FDF4CAB4C3;
localparam G12_5 = 512'h0682B773B8AA187AFD44AB4E6C4248CFF342F2FE2B06ACA6D7A05742B9CB855F1F98978D1D8AD412F4792106345FDC53FCFAEFE452A9260576C4A8DBF6DA3E60;
localparam G12_6 = 512'h00ABEFF76E8220834C463BCAA05B162E5001D9C73DC3F6F6250B4FFBE203591E043BADB0F04353907D24FE3A9F2E284F65F5134948314D8AA1E42C4A886ECC5C;
localparam G12_7 = 512'hC90CE07E4D5CF34ED33D18B985BAEAA93EB04BB6AE0A1EAB35E18791943EBC138666816489E609CED807BFBB040797CF761C1D56746956D5E6D1B2AF78F7D5C7;
localparam G12_8 = 512'hF5B7D5A79CE15C838D988A042755526D1FA555DD09422EC1F9DC1A0917C200E54450E8BE4F053ED4C317820462ECDF8F20F0B766621D24E41DB03088814D88A5;
localparam G13_1 = 512'hC0AF79257E31B3209F035206058DA1D026E4F6DF463E5CF19F6D222BEA741BDD09F9ADD088EEB7CB489E7BA21CACE4AEE1F597665AFAFF2F88DA50EB1B86452A;
localparam G13_2 = 512'h7EBFB2904CF9D7ECCBCD2CB98BDFA85F4F7A09597C5898D163B96D91DCFDB70BA03F7CBE46E505FF29855139DACBB4F2361816B7364109631BAB36AA71A7E560;
localparam G13_3 = 512'h2633191116F6EE689AC51275141A25312BB651D76F1A1423304BB84D51F07664846BC95C412B94208C9EA5864F1211B89D830A31168C866D68C1316D348B5329;
localparam G13_4 = 512'h93AB16F0563A448B474E2F1C30AC572B99AEEEF8EC13865969B09B30194D2AD9A45B77ACCA1F4586C7602802062BB450B4FCC6FF12D3D167709A5D48FDE85375;
localparam G13_5 = 512'h241C837190F9E8563885D601FEBACAC48F2D023DE91593196D3E54F52F661D3E29B67EF891B7AFC4121CE4E5B89852C6BE0EC09DC8B047ED18FB1D17E00874EB;
localparam G13_6 = 512'h0D0CE5CDD08DEA70EE3A7B207D1DF8D530B9ED49E7512BA69CAA0D72CC55EDABB138AF6B84F2CE4C247FF54AFD153FC1761889DC51FAEF5A948E165F8F9F8917;
localparam G13_7 = 512'h6C6807AF6BD56717C908E681153D715A90785DFDB9FDCB1FC502223A44BA29900F3AF2A56C9FACF5819EB89895220D517B3EE89678E04276EF5FE91CE0595713;
localparam G13_8 = 512'hC921D8DA283E0459E7830A45387CBA110608A45D5C7A44FF5656977CF199981A8D3C4ADC4CB8881B9E1659D937E16F3A3CA91F401C96279D3B1B5CA0630CEDED;
localparam G14_1 = 512'h7C22AD18A1E9BC4DCA2384DB32415770070F8E327F6EF485808D0ACF8CF2911ECC17D53A59D9602B26C6D39681855B5038E70F55DC5345E6D3DFAA2E97E70D8C;
localparam G14_2 = 512'h8933E2CF9E6D2698EC35523C8D03F5EFF3884E81859EA6A998E6BF0377B60855359E2CD955A518EB701E919A98222EF20BE7C4228AE933864CDF0F32A40F6CE3;
localparam G14_3 = 512'h398A0296F13659D46F8989D4C8FFE0E705F5DD862AC7C128C017A0CE1164E9B9B5E4768847420BEC856F2B060F00C083D138C12EC3CE2C2F3BF0BBB097B836FA;
localparam G14_4 = 512'h51B83E7F2B34DF0912B7C936C39E7EAF53323D1339D8B2B93DA1DFFBF051BF31C20DE9847BE9DA2AF41FFB29E07E87A29E4E2582900CE68B4E35C7D8C94924A2;
localparam G14_5 = 512'h738CA2519C451AB8C3D0EF773EA575D44F270F79A55ED6FE66460A28E0425130557F1D5AAE727BCB286FEE0ED7019EF97DDE49FAEDF022C92D29743AA7D01EF2;
localparam G14_6 = 512'h7C53289D362B97BBACA3A467951A8BAE693EB712A0B37648AF44F6ED8EC9742BA76D4CDC84D33934E1B173FE3A9C79129A12EC3E85B47C2410246EABEFAA041B;
localparam G14_7 = 512'hC62E5D7C354FB56F38C5D61B3C1E8CC96286CA18FBF79F3537A385DAF898EAE50DAA9593B8600179DFFB56195D419E81AB4F44739F962B2F85BA8C84889BEEB5;
localparam G14_8 = 512'hEC729C53D12F3630E3AA49CE1C93D2CA7ED03BAD77384EAAB1DFEED96F7797F24ED110BC0459E08518AB639ADC76DFB018C8841351544B8A47D9D6A132A057C0;
localparam G15_1 = 512'hF5E614C6079863817AC8472D454E43965D7BA90A2C323B17552F3C5916BC65DD3E84C5E4B9D0932F18BFD8D267473256FE1314497C08D81D854D84CDE05224A2;
localparam G15_2 = 512'hB4D16DAC333A447D9E00DED4B2B520A3F7C682A0CE1FD02514CBAF630E8C381BB468F86C1CE1485E8307F172AD9EBC0D788140A24F1282AD481F5AA2A7D38242;
localparam G15_3 = 512'hCBC6B0721996CB1CDAF70B76F63CA679308556DE592F22CFDB67C54E0EDE72C53D3698F9EAFC16EE91BEA2F6CFE450879020DD8551F607946BBF5991AA55DCE9;
localparam G15_4 = 512'hB377F2CDD7851A89A1252EEDFC05AF2EDBBB21F22696AE49993D946670F6F6FD1103D8093B39302A7424A7B923FA61BED6E71647FEF5E0F611548DB3992641D4;
localparam G15_5 = 512'h6FF2EE10D53B796369972FE29CA3CE81BDF62AAFBB66F517D0F84E9A92FAA3BA0780548035937D04CEB2866166784C2E0B34859E03D4CE4FF25C2E53BD86412D;
localparam G15_6 = 512'hA3F7ACC6F4FC9020AF5251B7872D9D6978E2A319C93BC311B3589C8C14DECA3B15DDA7E2D8EEA75B4125B7979F465DCDA31EF30A85222887600AF8635839E297;
localparam G15_7 = 512'hBF3D155E2AEE6E2099385FE1C829DCF426E8F476C7DAD3A1127F7765C5A92751967AF08498311065D1808823C7C3251D59A4B503AED60AFD2BD677D731B7C816;
localparam G15_8 = 512'h8BEFF5C4E7CFFCDBE0E5293B4DD5F925D40FF373E2FCB1260BB1BE5D1DF52936B2CD57D9E91F40E06EEFEF52A6A1623F03DE9A45325A324CBA058E111B3A6584;
localparam G16_1 = 512'hA21C8C26BA9700DD2A4C5A5DBE864A3A6C87F84CFC4D24EC4D799C78FDD33A4C6989984F5F94A6C83C322008111F95DF14A2B5121B5E5D0CE570A93E5EC5A6C1;
localparam G16_2 = 512'h536192D73B669D43DC0343C06E9197478FF62809CA7074CDDE873E9C9A8D962C4F9BAD702A84F1ED3BBEBF563E43CA231DFCA6D302A69DE6A78716829A5E4367;
localparam G16_3 = 512'h37EC873783774DA64AD75CBC81E7345668C82C1E4AB38D950833262FDC99F87707D9DF86B8A7FFBF10206E67261FE505A99E78DC99370EB4D6F439A0E369FE1E;
localparam G16_4 = 512'hF83FE12090AF478CB540DE88957FF008F24E0B3C9629871EB55A23AA1F18EE4CDFCEB2375EE26047FA726D13C2D08847F5C420CED73345B80A630C92C26F5CF9;
localparam G16_5 = 512'h34BA6D2C0FB21D7D0344D14E108B125DC8EF4BECA948D39836CC079DC4ED8FF2191F42397B1F1B58653BFA6319FACA6E2355952DF9255592AC97230411BFDDA8;
localparam G16_6 = 512'h00721EA63D1C09843A607BFCC8031E16D8AE2C876012A8DEA9C236B43B683D5AFB66407CB9BAB43755B06C746AAAD17539D332EEBAF0E5E2EB19FF477E8181E8;
localparam G16_7 = 512'h874E543A21447454EECA238420864865FCA5BE3002BF75DE1ADE2F5BF53AF506CBBAB92E76B4D54E637811261F244EA4631F57D69E13C5D43D167528381CC12C;
localparam G16_8 = 512'hC2F79544AB71014461F3181876418872E94C0FCBDD22331CC165F32A1E1090F599FF1E48BB2FE0CB5864F61A5B6FE81E5513617B7D7DA076BBA9692FFC6C611A;
localparam G17_1 = 512'h838BF3E846F3E52B3B1609B818E21D8AFE37B94914CB997B6D120955930642DCF847DB460D65CA6F70157CF5988FE6180146876FCDE094B34AC3EB44A9AC4BBD;
localparam G17_2 = 512'h8051D08739E2E5DA22250F01F6D09A92674FC918839B9FD49C1B2644D47F5FF552321B591C1A9595F96731F65634B2990F8443B72F3CB849F37B6AC79CC8A2BC;
localparam G17_3 = 512'h5118D99A12BBAA8A8E2A0AE50B48060AA22D76F57BF6D0D2658B7AEE648BF6F820C114933AE70D13F08F91561C4B91D355A1A8783648AB076931A7FCC4D1A92E;
localparam G17_4 = 512'h979C886D8591AE350CED09B9A78D8F6EDAD1E5D01BB261C244662BE4654B1E1263BCCBC78D62253A95C3BD6BEF46DF937DAAF2C1D3354D1742B0D3A49A96A610;
localparam G17_5 = 512'h8138678EFDDB6D70CD9F6166A6532B21E92E3367A05BFA95306DF0133488B1C70294022DBED7C46936609191F5944C85675CC09C8DB1B8036FF8CBEB53765A5D;
localparam G17_6 = 512'hE2E81231D905E55BA7D2D9B8FA725762AB2A3F67184874EF1FFFCD9BDFF2B44708818EC85AE2B30B6C82360258730CCDB229B975B35E8C8AAEF3BE0856E929A5;
localparam G17_7 = 512'h56594205AF5B8B62E8226F3248BF92417E9FEBC1A3EA192B2A724A70EFBA444C9F83612F503F6513B7088E5F0985388B8BE33A0A2F3E8883D08DDB45F8062983;
localparam G17_8 = 512'h94AB6C2A85ABAC52F23150271FAAA3C8308CE1AEAD42744FE6C1800F5AF065A35743AE87D5D1A4FF0EE3BAB43922106D9C205B9F6182F0B527FAB659640D2915;
localparam G18_1 = 512'hB847F4DADE720D0DF065DC1B3D18A7153D579D9A571C6EB4681D12857BEF926D72002B4E6F629E3C949E777D1452F941B24C2B6F84291F1FE16E418F55B727D1;
localparam G18_2 = 512'h11E84B7A3B6CA012D85B67D60780CC02A8D999FFDEB55C5481730F9E49EBC603968D88F99E97E799EC6E19757BE752C0E8EFFAC85ABF44B919BACF23584DE5DE;
localparam G18_3 = 512'hAC152E7123EE071DDEC6E4CF194C6CE9D0C9F50E083D44145FED3B039DD2DB61929DE81FF870CF38F0C476274D97DB04EDB9635C26464122C2137D478BECACCC;
localparam G18_4 = 512'h132173F581A4244E7D181B001C2E4C2B529F23F997D180F0B3E70E299D347B3B3120D4A3BE171656BAAF973FC6EFEFE569A21728F88573F0D977E62C7EBB221B;
localparam G18_5 = 512'hE6F13A94FF7142E1DCB00A91B10E4473ED5846A9673E2C0A4A0761536D2AF18FD0081A1DBB403255C14B3878E8EF4EBB256DE2CD78E87CBA6C2A8B7AEC6CA880;
localparam G18_6 = 512'hAE6308C2B679C77B1CD3032DDA4D4A6C07EE83A3361EDF53E28E5D300F7E2FEEE2BB2B92C596179699D8CC2166F30E602D47468781E691B423D6A4E81F19C11E;
localparam G18_7 = 512'hFE685C3C6253DA415E9AB859380BFE7F06024F31CE177BC9613561F7900682A9DEDEB41E077AB5032878CAD22F3D41309E1E9FECA8B91A331D316DBE7DC40534;
localparam G18_8 = 512'hCDD8754E6914EA86370EA93B19CDDCB0E73F4047E7875FFAFED8CF9F4B0EB10110DC3CC90B1FC74FD90917760B616AF08766F9C91C67E38A81FF05269A937525;
localparam G19_1 = 512'h47C094E714143DE5742BEE47211454AB3831F336409EBAF1B0758F406742353F2398C9EDA2B4254E791485A4D42A84E18E959450121440782B0FBCEEDAD5FCA1;
localparam G19_2 = 512'hA434E3A99E4FD9CF2CE721D66FB7D42034AF237A1EECF2092DF066A1C55526749D2E328F0C556DF4FAA503A32CF9558BB7F85119168DD421B82C21D35DAD8986;
localparam G19_3 = 512'hF8B39F5147B292CE7BBA0D00B7AC51053B5E88DC1280348CC3C1A173AA113EB50A6BA95E0E7830DCC91EB404A3A11C74D4109D8F48AAF575A57A86005E38C0E3;
localparam G19_4 = 512'hCF084E76C7E361F7BBD9E38830649AB6795246C810092A8E251191CFFEEFE7E87FF0BA2D77290349E77A00E0BAF1C30C947EC7AE034A97A094941BB032BE1A7A;
localparam G19_5 = 512'h29DA9C1A2C41943FA65425134FC926DA62192E1C692DF3A0F3E063EB282F91A1A49DF5D0B3AAEC8E5AC8B7BFFF2053279FA0AE563B0186701D8A57D325016CC6;
localparam G19_6 = 512'hDE1AC50539874615DFAFD011CF7227060CCB69F13BA8E128B7A82B33704A5C8785D359654D31242A36A9EB335E9A595E925BA288181F24AEE09F40F4D9905964;
localparam G19_7 = 512'hD88D0B9555FB77349DB1C44F3E5C85F0ACCCC7FCF115B298D9914219B253074610691D9D28866E107D1F84EEC34E692CD0E2050B60C6D193040D21439EAA93C0;
localparam G19_8 = 512'h0E113B8B6EC30804FEFE51792167EA29143D3092FAC3C1234F4AAB57CAFB4A82AC0C20B3F1EB3AA32FC7F4B07F89DF965375614A4E0B013EB362E3FFF7064841;
localparam G20_1 = 512'h70FFB209619E4EFE3FA9DD7178FE4DECA4C6EB753FBF191DDE03F16F887BC9782DD4A13B06A164D27F3D1AD92698EDD78C6392D340FE1E68B2069CE3F5A5D77A;
localparam G20_2 = 512'hA2037223BEEC4F438F386721D814DEE5C121E76F1FD638765FB1F1286D00AF73FB22D84E71816663A61C50B77CD4E4F6208ABBF6ED8204F874EAF2C7183C7B37;
localparam G20_3 = 512'hCBDE288B44FF3B1314AFFE2708D04D80B877E93CF1B7A2ED64AFCB38BADFE6732EFDF24A88DEEBEE8A47F4827483CC3A60AE6C41C0EDC33A004B1E29B62865CF;
localparam G20_4 = 512'hA1DD06F5F1B6DE558271052B1239F171D2B6BF58786560C83A620D7F6531C4FF94AA82E5FCA00D10FCCE1C74358ED92D4D9A6F3BE04B6176208112838572650A;
localparam G20_5 = 512'h408A4B428C92B387D75534AE21744CC3C30DB5C97075608292713F68B6814E04B3D976055BC90B40639B6950831EE910D9D5414F5BD79E05394D50B8D2E7410E;
localparam G20_6 = 512'h8E8F06B7B76F6FBB52C12DCF274E9438727577356E3D983BCA4E2E91FA6E6EE26D07E7FE758CD2293A92B0466CFFC8A972FE2D51361B4CABFF3B2F853FD0466F;
localparam G20_7 = 512'hCE0CD09FC1A9E4FFD6E9898951CD8F354CBB12A08550E5294A45E01BE01D965AD539CA9EC5912C890751A454169E1C089B06A94E3B5F43CC9A189626ACD3191F;
localparam G20_8 = 512'h980226CBF2CA0E8DEB4967B70BBB329194CC8DB14AF9970C87BC5FDF246BA31CD30D4515E2D65295EE08B86886D260E14F93827A7A8EBC347EA8AAF45ADCBC9A;
localparam G21_1 = 512'h43DE7A224F0FECB0FBF13E3D73F842BDF8C721BE5A03406FAF104E3CC358CC4533346904671AE05D5E724DFF08CD5D52CD22C1A8E6778390CC5FA783D096A193;
localparam G21_2 = 512'h77D7FAE7B12DE8CBA98F1BDB3507B52033A6B0F93C0B3435B3D57220606A04F3E09EB26E98C5A71D636829623DD9026B1D86F0DCBAFB091A030214583B8B1B0F;
localparam G21_3 = 512'h5A8B748DAA524BCE91822B77E9913A79912A4E275E3F891153F854AC896FC044FCECBAE7557E67781D9CF2E3C05054FB052DB366B94828045616BE3C8A60827F;
localparam G21_4 = 512'hD13FB7359642A94B48DB9E9BB5A69465EC5737C654BF3F13D589E7C41894EB7C92BF3A4C770163367552778CF13E8FD17A09363FCF67F70FC55BB53406461891;
localparam G21_5 = 512'h076B6655C01A6A9221887A4EEB0022488F572FED49BDAD1C02996163B904B24C6BE4626EA82532930768EC5241CAB37098C83EFCA76B6E753AAD3DB45944BDD5;
localparam G21_6 = 512'hDC4699E4FB1A6F5A461051395951E2F807761DF909D92C842E481BF9DB1DEFCA11513B1B379F1B96281DDC65644756A54907567F280F3D5D7A9681C5B48594FD;
localparam G21_7 = 512'h1665DB277BB3619BDE1237C37B02D4EA00AB22E7904AE7C4611CC57C5AD2C12C358968FD8069B3D0F37D629013F0E5376B9C46E2F719291B4229005F15C8BF55;
localparam G21_8 = 512'h3DEF03EC009E21705ADD10B220423367D239E13007FB20D9DC7BAC093A06F949D66E619C141DD265BE0D807EF86F2E36C16690B5CBCBFAFBC3895BC80DC6C717;
localparam G22_1 = 512'h2FE7CF36F03952549ADC923D606E8B8B75F6AB93C3E564F54E21B702870BFF6905CFE5231E6DDA794BE56D45779E808E88346F8DAC3F08A51E0197C088E4F541;
localparam G22_2 = 512'hDF4B156899E2068C4ECFFCD950C1B1B0BB7D2D382D03578DF029743A1D22D7B8579C2446650CDBC8C3438EAC744718B70A00A7616367570A936EC8A34295D432;
localparam G22_3 = 512'hF9D84A4E2E6EFFCA516C3835C45B51091C77DBDAE5706A57A3EE600BA423128C33ED75E1F9F2CE7FADB85EAB1F8F798F320C9A322EFC1F5DDF2991599060A64D;
localparam G22_4 = 512'h57CAB93C1A6B3B73E58A9E9008C3543E01294C4CB491D62437466DA61263DCE085D40C6C19EACBE95D92850751BFF88BAE4BAF74D365C85D29EE0CAB53FA32CC;
localparam G22_5 = 512'hEC617100FFF4AEEEF35E0628C82A5861196003C7BCF0ED7D6E747A7D2980F292A208FC4D7DB8F17CD9082891167CEDD28D9A7A1A50AFD382C8C77F1515721DEC;
localparam G22_6 = 512'h34F9DBD9A9F89B436E63C7D1202F2D83CE0EEBB6C1FEE18F4EFE838278F54F5F8CEC9C8183C1BA03E94A554B2B6D71B70673DA9249ECE7D7D3F1ADD0DAC7BC31;
localparam G22_7 = 512'hC8A01BC7F86428C6EB7A2A06ED49B50B7D0FB253311D01D7DD77445F29E947AA3E9D9DFB27B10D7E532C9C56E19C63068DA7BAD03284C486006DF990B72696E3;
localparam G22_8 = 512'h7BBBB5626C0AF1DA12C7F8955D2A9544E5E85D51FE4F0CFF808CC147493DBC378D9A1AEE7C8DD96E7AF78375AA5AD1019CF892C9E13586F6722612A70677CD4A;
localparam G23_1 = 512'hB5FD20CC39FC444C5F72C506C41B34873B588321BA720FE4A157C8CB0B3DA464AF930205ECB56C458E4C51AA96103F9A9C393C05437ABC4BBD4D7CC801B0B12D;
localparam G23_2 = 512'h03B90C3C218B63FCBF5BE95352BC90A75112661622A2B820239D2FA0AD251173D9D4035AF3DDDBEE862A46E4E6148C7C07C4A9BCB843672845B9C971AC2E0627;
localparam G23_3 = 512'h1AD2D5B81178299D15D4A05F62732A1512403C24DA7D44067807705889A0B746296BB7D6331EF209E28F23BB89C8CA6F76C25ACDDD8DD663AE8F8BA59B7A473B;
localparam G23_4 = 512'h7F9396696A8CB753C8B50CD407D90C3FEB6C777358DE22E926CB56660710065F065B792342EFC8EB4668EE4D994E96CD8E19D5FAB19C8AD6734DDD3E3E06C64B;
localparam G23_5 = 512'h721D4A6CC537BF3B3FB317BF9DAD31E65040B8324D1C8C8252D144CBAB2F1EE8B3D1E8ED1EEA0E4855EFA4912559C2F48F563537FD2B0FD5ACC7EC47CD0E3FEA;
localparam G23_6 = 512'h55E6A59CE67BF6E649675ECE3442FE63BE4213390B886363647F5380A282E71F0D7E84342AA15B318C16615F6F2AACD2D3F5968FA945B194375EC4D6DF37DE47;
localparam G23_7 = 512'h40181281BF74696787C5AAA24BC4D456DD34550D70AB856004DE793E2745C5186CE2FBE7483E258B099913AC2145284FF1130BA07146A4BDB198FD48CAA76862;
localparam G23_8 = 512'h7C729D639CDBB755DC1742DCD042518689AF31A6C5EAFD0AD24425F2D6B42D29E7E0C3CB2EA2FDD188DC87AA4630AABB87449A093021455C99D9CC06FD413905;
localparam G24_1 = 512'h9CC642A176B98677B7DD6D95A688AE77A0B6CF3815CFCD4418CFCBC2981167EC98EA5814E8C4C0C4D82F9E22B2F234E3A5B33FF0E015569F961E1BDD5FB59E47;
localparam G24_2 = 512'h57492BEAA182A05C5BBDD8A04E30ACBE6CB8C04781ADD43E0A90296836FFE1E3391EF6FA38FAB30B49DD4BF00875A670D041557FCCD7F05706045D5A7E923EC6;
localparam G24_3 = 512'h256422331BF3C0112C4E5DBCAD76B212ED29EFC33D9AA553ECC9F8D138E3230D5B4B2A46223DEA20DBC9D86D54ACC75144BA528DC45DE611EFB5C97DA484FAE0;
localparam G24_4 = 512'hAEA86017E52C60A576BA4352062DAB7AEC292EE3115C72D7EEE62FB2119DE7B9E8BE01802C7DF16B0AE59566A75FE4ACEBE44ED7A36ECCC26499D000E8AA3546;
localparam G24_5 = 512'h2764DF6D7BC61CF7E9DBB65260806BCE27C647E18764C6BC048F7C0EFD14415A1DF3E4566740866AEEAF3731D31CB6028B0395E88575BCF3636D3437899A8A46;
localparam G24_6 = 512'hEE0073E2CA1BC867B02B105E6F17C2A41E5EC56BCC1D0513E17664FD392EDD1E26FD792280344E03CE7BC758EFB37F785627E486714182B4E1C16F103F892107;
localparam G24_7 = 512'hAE287A4D57A3DDE70DF2BF6FD30727A7F5C4256FC69D075F3895DB2B7C3DA9BDB4A082A409B466549AE8BF39DEB7516D2712F6C912423A64FD8A3EE50AB1925D;
localparam G24_8 = 512'h6CB58E5D9EDA695AABD5989FAA6F0E6BE69F4E6D843349CF509FC9CE8AF9BC39C54079800DF7189FE759FF7623174DAF06049DD4928456BC9D5A757224B2096F;
localparam G25_1 = 512'h616DB583006DB99954780CD6DFC9908772D8260D390B1D462A8F62DE8809216194BE0531EE408AEAF27F50F3AD71865AC7910EEF8824A858CA7B13FC843DAFB1;
localparam G25_2 = 512'hBA3E0B010860D09066A8632E2B273DABDF90C26FCDD989C2831874EA7FBA23D940A294111C1B0C1CF62F56A376B94CF64FA594B987B19226E525704D7F2BC66E;
localparam G25_3 = 512'h226C671C22A59AC062490596EB1536C9F66AE799C2489FAD2C131E29ED64A25CB0ADC88D04C5EC8FECD7F78B3825E626858CFAA0DE77772CE8822C7AA39628A0;
localparam G25_4 = 512'h123B1C426E2A93366D067D26DE51362EA0BA916EBD1229521B1B044459B325785F3F3E24199B2460151E4CAA9FD26A5DC46BE0D6DA907EFAF38F413642F702F5;
localparam G25_5 = 512'h324AFD5D62F4CC251FF5C0FD95DE0FAB061F0C92CA5BC97F976118AD84E0663A3BF1B4F07D1CCCC2DF9E09D506B073DED87CC0653C944FC7D438223C0DF3EB67;
localparam G25_6 = 512'hE62AE13F8D4000D616E814045495F6E969C473B059386F5DDBCC25F4002EB132D73A98414D85346F55DEBFF875F7CB9D2466A412D180E0A1ADA18D281376A671;
localparam G25_7 = 512'h8EB0FB6BB7B9AD2A2132010511077F6BD424B6F5B578C11D0076B781930F755EBB72C41ED17519476C257C31C3159BF31FADA2755F1B8A23B22D6A428AA290E2;
localparam G25_8 = 512'h54CC73C7599AB67C6807C4286BECF8423F3216EF04E1B6DE61349DDB23E3A0EB0EF70C5BE1AD91D31B0BB532C1098DC619BF80F3853EEA357091C05D95170A7E;
localparam G26_1 = 512'h5E6381A718C0A817F8101ECDCDBF825E732E4356CEC42C222DBC476BD704837C382B7FBF282B739EDC22B5EEA2909F0EB3ACB9E41FE2AC791130A36A9CBFC1D9;
localparam G26_2 = 512'hD4F8DE28FA77F37E4A6B5A82A58CE917CA74C8397E9DB8EDCB2BF65DB91954457707FE876DFF812D4B99466DF479A00114F27E702249DB3E9311301E9CE98703;
localparam G26_3 = 512'h74FEAD0013FD861D67D7CE69D3635ECC6266E862D08B63077B45D3098306EA74159DAEA2263E58705EA5ABE58B7FD41862B9EC1D0F1BD47CD6CB42739C24F7FE;
localparam G26_4 = 512'h7ACFF6D64C8E8F94BEABE280CFDCFCFB26AC7330073C25E0313DCB75E6C5261F15D82AFA665F73A4B4DA4E5D1648EAB051EDEB9857C13C2F019FCBBA4F9DF2E1;
localparam G26_5 = 512'h9CEFF1147D792C14AA2E211C3B9B94B2C9F24F49B0B1ED6E200C88D743F5AC1EE283C3A0AC79B9F1F496BDE74A2AA591ACF2F526FB24413A58B495F91905F596;
localparam G26_6 = 512'hD8F1469BCA9CC5041C50F1FB479CF2680503AD85BA2C0C6D01D2D739F3129315E49A9F57236D9585CC0B8A9B4BFE9ADCD97BED9006C33976ACC00468693D56FA;
localparam G26_7 = 512'h1EE66371B0EA6C4E1E172C2C5D76806CB7376B8CDEAD96B14A1EC2B656298B9425EA2F0671082D70AA23C267D1F215C59239AEB40186DF0AB284625DC6BAF45E;
localparam G26_8 = 512'hFBFBE26BED98BB3B697764A6F82C94039CBF14CB538A7D87801ACBD3A444A858BB74F0A4707592EE6B7DC6D21B8F6B4A184B567C8AA4CD825EBF7F1EDCE015A5;
localparam G27_1 = 512'h25453670647D23C5E445A705953F3BF4A5AF02E7BC46C969C8141D8782F171C9CFF7EBB20945DE5D363AD36D3BD5A0BA081C079CDD04B6E5968187C8A665344A;
localparam G27_2 = 512'h23E9B1897A6FDF427B5E910AA8D71F9CC6351474BC4563C20FD38953295D3BA15E7D1010503B7BA1C148251DB8A88AC64E6AF8C1CC056E4EEF1C927FEC40C35D;
localparam G27_3 = 512'h57140969483D9E33429FAFD177D031A43B727CF832C8DFFE8D8960CB55BE4BE27B69CC26F2FB731B53250D6F8EE7DFDA98812B9AAE9C02AE2FEDEA598D6B6E2F;
localparam G27_4 = 512'h22B6CCA50541BD9F5D48565E551B310E10A0DFCB8035A5EC86EB9CD8C811CDCBCCCEC3732EF93EE8C9418E25CA5744E07C45F9B161E277BCECE388B9B84AAEC4;
localparam G27_5 = 512'hDA37FE277C72CB5CB1BE92AD373867403E46B3535159687ADC79C39DEF7005C1F11F1CBD5F8877DA66AAC156EF27BB893F5F1132336D52E8AEB60EACF9BEB3CF;
localparam G27_6 = 512'hD204D92DFA496DAF564272E3FEC51CE53C8F2DF6ACB191E60E14CDEA28FD5ED0EBE09672ED11A3F6466FE3A967A4EC8390303059AE00DD83102A9F33B2943E4E;
localparam G27_7 = 512'h6E56928E7FEE3333A36FF3EE7598744CF7C298FEF3EACC7CCC0F36DCBA6D87BDD441081163A65E27C958AF79C33A98B81814015E77F82EF5120FBDAB540893B4;
localparam G27_8 = 512'h7BEB68CC37F23835C91F5D36D6BA6F0A5E68FEBB6E6A2F247EB5CF57684D0770249460788DFDC4A1218652BF881B4BB06308EF86484E7070AACC72D3977CF5D0;
localparam G28_1 = 512'h6230DEF1ACD4425F7B155A2A285CB2A32CB9D46DA09B28167826E77AEBD85F0C416595E136184841451F5B3E1F17D02C3DB32C2AF50091D6376406D8CB78A9E3;
localparam G28_2 = 512'hD3B19911ACC450679EAE25B0F290FF372300F1A4BC91A43CB79DB270133D41DC4970F1420E71C0F816EF938C3C17F0FCBB6E920ED853EAF6D2DC6792BF87098A;
localparam G28_3 = 512'hB94C2E5DDE78C974AD6F423CD5ACA01EC9420AAF3FE83BEC31D47AACD3D62FA2476C38595BD66639368181E75B44BAA7ADBC2B42E1D82D7A59312BB9A16F7D35;
localparam G28_4 = 512'h0B13B44D828071E69DD90DCD9B713A05FD8C21AA5E6E6D8DA49A5C3B34F98A4E5E822513F0DA200235C65BFCA1DC2CE4AB21D146B778F6806680B8AC75285760;
localparam G28_5 = 512'hFEF66B861AA67C768A76D585DFADC8EB6556AD841DEA9F44ACB42B6016142B6B69F1833474FADEB0400CE4D9F3BD62AD96E57F3E93DD229180F2D4B5E77D098F;
localparam G28_6 = 512'hEEBE2DFA4D4D86ECB07EEE9565FB589855E1F53BA1B9784A8D195A0E3721551270089C535216636FBEB4D9E50A9EAC3DCB27891A7005A2AD87427E6B8326F6B3;
localparam G28_7 = 512'hCA225C7B2A9EABFFDDDBC130B5342917848B029917BA98FFD6EF2389006A6B417F678C61458EF625C96C0D3D07945ABB9836CF80823EB6244D86D114CC5DC2B1;
localparam G28_8 = 512'h94F5D55C398B16A71497C4CF102C2F1035C19D5DFC8A301B8DE33D41D909C15A3093B09E7489CE6AA14B331B70E76637FE6DDFFFA6DC4C510371CB0D2A6EA3DA;
localparam G29_1 = 512'hAC5F866DD75CD4C2D5959AC37DE4E1E870313A5B2902F234CD939FE39F31FEBF8B46DAC906E3EBA9C3A74DE46E7A9140D3716667BB1EC22A87D5F8D048BDC5BA;
localparam G29_2 = 512'h57B6024327CDDFF3296BE6508C48045B71FA519156F8C125F4E3B7356576F32C63BC588908C4E8B3F9F2D12A9E8F35B6FCF296C17FD8E8D076406FA11D16175F;
localparam G29_3 = 512'hCC45AE82D672979E8A0A359B2328C79AE61F87EBE04DAC9343030548659732000CE627417B3F8CFD4A992E7F2B680216AF773385B9337E1743D43FD965282CF5;
localparam G29_4 = 512'hAE71B0CAFEB4DA3E0B95F1341667C519FB9F89D7CEC711E57485F04A965CDC832CBEC0BE1B2A3E23B5EAF4C5DAD8767E054B2225A60B88BE1DB6A35E0BAEB237;
localparam G29_5 = 512'hA206BC721B252D52EA1F8E311203DFF0AE8D65BD1986055701A3C7FEB2DDEDD2D57C3BBA6A2BC56A9157677D7B48AD2907927176F6B22E8A92F6E9863C9E16D9;
localparam G29_6 = 512'h11B6209E06EFE6ACBBBA2214EF5AEAB9D76645476B2C16B8D14E1AE3F3A85188835922B914D3F32FE05B7987A2516B3D3C8983AE176DFD04349A45359B422E1E;
localparam G29_7 = 512'h01CC2266F2B68A4323F8931D7AA37B1CBD70DC2FEE91592327207AA6121795150A0DC918704A1A293778FE75A99FDCE77E820D0905EF7AC72A682F2487A6E0FE;
localparam G29_8 = 512'h03F42D94FDE1C13F958DF61112DB4A27A8A8EF35087FD089729F0864C2706CCB2B6CBD91A9A7B7B31E08EA3570A6E1BED495FC84FACD829F3234B1D1DC574B67;
localparam G30_1 = 512'h900AA496432959141795C615CBAEA98002440A0D447EF990435E452CC690203BDEBCBA3EEFC7A7CE71EB54B1728AEA9EDE70A7E6A1A8AE86168709A899738CCB;
localparam G30_2 = 512'hC5B7A094AEBEA8EC95A414A8DE5D3DBE6745CB0D330B78435AC2BB6666BB2D43A19EAD3B3D9536D0BB92DB949570981C22805E7DEA452FA649C84EDC4324A7FB;
localparam G30_3 = 512'hE6A9CAF4EE48400720B8F84CAC3A42483B7E571846E2A5F77A983EE311179CEC2D99878FF5AA06ACA0CBBA63B36985E0970761E7F837650BC46C9A2EB1AEFA95;
localparam G30_4 = 512'hAC4D8AA5C970BB55FDF3408356C9EB2683B6FEE593736B66B49C055BD6503EEF3C7CADD15C9B86DCA626E1ABF4B971D04C0A9A5AEF8305C3D0E4CC02C32FA91E;
localparam G30_5 = 512'hD8949EF8FEADF7DA39D395B52D2779A0B305C4FD10C33A434878967D9321B4835C035CA5802C37F6DC1E39AC30337253114176BBB26576317C72E9548F179A5A;
localparam G30_6 = 512'hA200FC35B6A0934D57543A60F6114B7B0D78D8DD8932538E545D806A1D9E47390F092501F4A470CF7B1F9144D0A8F1B0C3D607930A75E5A150233DCEEDB4C10B;
localparam G30_7 = 512'h217C8EB38D4D2A0EF12557321D504ECA670B41E496441FDE341F0232101D4E3F4158FF6F4EAECC073AA811DD450F528BC6095868B7BF953926056BD409E5FE36;
localparam G30_8 = 512'hB82831B150B80A736D6CF7B16660ADCD5E1F4DB96E36E33DCC2F1506C7B8B0F2A4EC362FB0CF7B8B3B08D6CD1AF7440729D4C3C02627AD8733A0C94B2EBAF526;
localparam G31_1 = 512'hFDB4463E6F8FBAF565B1C3320F5704A87309E529842378ECB733784F1CBD85F4F87FB0525C7C4D307061F74DE2FB3BDFBC77E04EAB75A64FFE51203AB925E807;
localparam G31_2 = 512'h1D1101A16A2C41DBDCA94C128560BEFDA4ECA6F22B44C6E5085A23F84106E4FD870FAA789E03FC37086E67B69FC8EB6421AA57FBA27866DFF712D5FEDA21FC51;
localparam G31_3 = 512'h76EE3CB2C4A8629C20FC646A7ADF2A4BE73DCEF53FC926067EB9964996BCEE403C5642CD2F8084E0C14D3627FAD9F0180DADF07331246C007F3AF95CC9B451CC;
localparam G31_4 = 512'h3638887EB493F5EE3361F07E00F115BC04AF404BE6BA3467322B37A8E6ABF47710D56C3BC751892CFD12F29CC4319D0562005562D05261D39FDF528A11E65BBE;
localparam G31_5 = 512'hA0BF07C52E9A9ED7AC3F0FB9196A450E162009509F20BEE74FCC6316BC4824D93CBAC25E470A7468A629EB520E980DE31F8C8873F4ED21B57AAEBF43A5754359;
localparam G31_6 = 512'hCD089ABE548975678C2123223CF3F345AE0CECF0A3726BFBB130E34169A874B6C4CDEFC0A05D7DA1EE475E5407F1535399086700874C13000E2EE21DF3EEFB65;
localparam G31_7 = 512'h4BEF6F2B4137DC6EF197D514E904B8F31BAD6C846D6BD7D7480F4818C3C57B4C7F53F168E48020273702071EE48EC53422C71C90AA0262982B82BB6FF3100D8A;
localparam G31_8 = 512'hEB3E8F033DA73FA82B3B93E50C60E5936A07D3218946588D0EFB39E1A55C0FB9DBA87DA50C4697EE2ED72B004301019E595B92A2F55F7F1B37C2030B79057F52;
localparam G32_1 = 512'h59CA13359E16B10A7F8778BBAF5D45E32C643B524022FE777A8F557C14141D638E84BC4DBB1CE5866CD0B89C1CC5C6F7BF7E25D2B4FC28A16E67CF8BFAC4F4BD;
localparam G32_2 = 512'hA612F30067700487B6584B1AD578659FC2B7443228B2B7B443882DABBF55739CB9660F530631A2CFDCBE94D21692CAC01DA9EB5048FFF17BC4FB5957E8C9DF1F;
localparam G32_3 = 512'h29E0573D85359FB7924AABBDDDCD26F5740FFA6824FCFCBD53BF1DFB587E0667641DD3F82962F5E6EA26461279B0F69479645462983DBBBCC544DA90255121EA;
localparam G32_4 = 512'hA97C7B71923F0382DF60C9E34D84CAC289B578899EBCF924F4304B80581C9887B1198F074143DCC4324D7DF301466AC97903E688DD2E9186EDD2D90C34202AA3;
localparam G32_5 = 512'h90815D489B715FF604788F335322DF5C8856FD85F753785A96F4B2561990F458C69D3F99A8ED1BE99C3F5A14B19B37AC729B3F35ABF52006E814B597145FA3FD;
localparam G32_6 = 512'h86A5A2038BB67CF8225BCCF7A587E0D09B47D26BC4DB017F6A77B6DEC5AF5B117E399D8A336358D4AABE9C8E7EAAF6447638F2DC66EF65C100D06EE202013042;
localparam G32_7 = 512'hAD845A43D23E66FBA72D9D56457D66C7E44D98ED1E5F1D063A5D01043930E9C2EDED8BA9DEE5F9DFF91CD887F097B9A2DF0099E278C253E0A549C7A2D81078C6;
localparam G32_8 = 512'h680566EA7A1E724A99B5D7099AED278A3065BBC64BED441154DCD346D38C9771648D55656B16CF012D0C6EC8F616D3B758089A8147D731AE077D557204256F93;
/***********************************************************************************************************/
input clk;                             /*系统时钟*/
input rst_n;                           /*低电平异步复位信号*/

input [width-1:0] s_axis_tdata;        /*输入数据*/
input s_axis_tvalid;                   /*输入数据有效标志,高电平有效*/
output reg s_axis_tready;              /*向上游模块发送读请求或读确认信号,高电平有效*/

output reg [width-1:0] m_axis_tdata;   /*输出数据*/
output reg m_axis_tvalid;              /*输出数据有效标志,高电平有效*/
output reg m_axis_tlast;               /*码块结束标志位，每完成一个LDPC码块的输出拉高一次*/
input m_axis_tready;                   /*下游模块传来的读请求或读确认信号,高电平有效*/



/************************************************进行LDPC编码************************************************/
localparam STATE_waiting_valid=4'b1000;  /*等待valid信号*/
localparam STATE_data_out=4'b0100;       /*输出信息位*/
localparam STATE_waiting_ready=4'b0010;  /*等待ready信号*/
localparam STATE_check_out=4'b0001;      /*输出校验位*/

reg [3:0] state;               /*状态机*/
reg [$clog2(n):0] in_out_cnt;  /*输入/输出计数器*/
reg [n-k-1:0] g;               /*生成矩阵当前所在行*/
reg [n-k-1:0] check;           /*校验位*/
reg [width-1:0] s_tdata_reg;   /*输入寄存器*/
reg reg_flag;                  /*指示输入寄存器内是否有数据*/

wire [n-k-1:0] check_sub [width-1:0];
wire [n-k-1:0] check_reg;

assign check_sub[width-1]=m_axis_tdata[width-1]?g:0;
genvar i;
generate
for(i=0;i<=width-2;i=i+1)
begin
  assign check_sub[i]=m_axis_tdata[i]?({{g[sub_size*7+width-1-i-1:sub_size*7],g[sub_size*8-1:sub_size*7+width-1-i]},
                                        {g[sub_size*6+width-1-i-1:sub_size*6],g[sub_size*7-1:sub_size*6+width-1-i]},
                                        {g[sub_size*5+width-1-i-1:sub_size*5],g[sub_size*6-1:sub_size*5+width-1-i]},
                                        {g[sub_size*4+width-1-i-1:sub_size*4],g[sub_size*5-1:sub_size*4+width-1-i]},
                                        {g[sub_size*3+width-1-i-1:sub_size*3],g[sub_size*4-1:sub_size*3+width-1-i]},
                                        {g[sub_size*2+width-1-i-1:sub_size*2],g[sub_size*3-1:sub_size*2+width-1-i]},
                                        {g[sub_size*1+width-1-i-1:sub_size*1],g[sub_size*2-1:sub_size*1+width-1-i]},
                                        {g[sub_size*0+width-1-i-1:sub_size*0],g[sub_size*1-1:sub_size*0+width-1-i]}}):0;
end
endgenerate

generate
if(width==1)
  assign check_reg=check_sub[0];
else if(width==2)
  assign check_reg=check_sub[0]^check_sub[1];
else if(width==4)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3];
else if(width==8)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7];
else if(width==16)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15];
else if(width==32)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15]^check_sub[16]^check_sub[17]^check_sub[18]^check_sub[19]^check_sub[20]^check_sub[21]^check_sub[22]^check_sub[23]^check_sub[24]^check_sub[25]^check_sub[26]^check_sub[27]^check_sub[28]^check_sub[29]^check_sub[30]^check_sub[31];
else
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15]^check_sub[16]^check_sub[17]^check_sub[18]^check_sub[19]^check_sub[20]^check_sub[21]^check_sub[22]^check_sub[23]^check_sub[24]^check_sub[25]^check_sub[26]^check_sub[27]^check_sub[28]^check_sub[29]^check_sub[30]^check_sub[31]^check_sub[32]^check_sub[33]^check_sub[34]^check_sub[35]^check_sub[36]^check_sub[37]^check_sub[38]^check_sub[39]^check_sub[40]^check_sub[41]^check_sub[42]^check_sub[43]^check_sub[44]^check_sub[45]^check_sub[46]^check_sub[47]^check_sub[48]^check_sub[49]^check_sub[50]^check_sub[51]^check_sub[52]^check_sub[53]^check_sub[54]^check_sub[55]^check_sub[56]^check_sub[57]^check_sub[58]^check_sub[59]^check_sub[60]^check_sub[61]^check_sub[62]^check_sub[63];
endgenerate

always@(posedge clk or negedge rst_n)
begin
  if(!rst_n)
    begin
      in_out_cnt<=0;
      g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
      check<=0;
      s_axis_tready<=0;
      s_tdata_reg<=0;
      reg_flag<=0;
      m_axis_tdata<=0;
      m_axis_tvalid<=0;
      m_axis_tlast<=0;
      state<=STATE_waiting_valid;
    end
  else
    begin
      case(state)
        STATE_waiting_valid : begin
                                s_axis_tready<=1;
                                if(s_axis_tready&&s_axis_tvalid) /*等待valid信号输入*/
                                  begin
                                    m_axis_tdata<=s_axis_tdata;
                                    m_axis_tvalid<=1;
                                    state<=STATE_data_out;
                                  end
                              end

        STATE_data_out : begin
                           if(m_axis_tready&&m_axis_tvalid)
                             begin
                               check<=check^check_reg; /*计算校验位*/
                               if(in_out_cnt==k-width) /*本码块的信息位输出完成*/
                                 begin
                                   in_out_cnt<=0;
                                   s_axis_tready<=0;
                                   m_axis_tdata<=m_axis_tdata;
                                   m_axis_tvalid<=0;
                                   state<=STATE_check_out;
                                   if(s_axis_tready&&s_axis_tvalid) /*输出本次信息位后,需继续输出校验位;若输入端具备有效数据,则将有效数据寄存*/
                                     begin
                                       s_tdata_reg<=s_axis_tdata;
                                       reg_flag<=1;
                                     end
                                 end
                               else
                                 begin
                                   in_out_cnt<=in_out_cnt+width;
                                   if(s_axis_tready&&s_axis_tvalid) /*输出本次信息位后,若输入端具备有效数据,则将有效数据输出*/
                                     begin
                                       m_axis_tdata<=s_axis_tdata;
                                       m_axis_tvalid<=1;
                                       state<=STATE_data_out;
                                     end
                                   else
                                     begin
                                       m_axis_tdata<=m_axis_tdata;
                                       m_axis_tvalid<=0;
                                       state<=STATE_waiting_valid;
                                     end
                                 end
                               case(in_out_cnt)
                                 sub_size*1-width : g<={G2_1,G2_2,G2_3,G2_4,G2_5,G2_6,G2_7,G2_8};
                                 sub_size*2-width : g<={G3_1,G3_2,G3_3,G3_4,G3_5,G3_6,G3_7,G3_8};
                                 sub_size*3-width : g<={G4_1,G4_2,G4_3,G4_4,G4_5,G4_6,G4_7,G4_8};
                                 sub_size*4-width : g<={G5_1,G5_2,G5_3,G5_4,G5_5,G5_6,G5_7,G5_8};
                                 sub_size*5-width : g<={G6_1,G6_2,G6_3,G6_4,G6_5,G6_6,G6_7,G6_8};
                                 sub_size*6-width : g<={G7_1,G7_2,G7_3,G7_4,G7_5,G7_6,G7_7,G7_8};
                                 sub_size*7-width : g<={G8_1,G8_2,G8_3,G8_4,G8_5,G8_6,G8_7,G8_8};
                                 sub_size*8-width : g<={G9_1,G9_2,G9_3,G9_4,G9_5,G9_6,G9_7,G9_8};
                                 sub_size*9-width : g<={G10_1,G10_2,G10_3,G10_4,G10_5,G10_6,G10_7,G10_8};
                                 sub_size*10-width: g<={G11_1,G11_2,G11_3,G11_4,G11_5,G11_6,G11_7,G11_8};
                                 sub_size*11-width: g<={G12_1,G12_2,G12_3,G12_4,G12_5,G12_6,G12_7,G12_8};
                                 sub_size*12-width: g<={G13_1,G13_2,G13_3,G13_4,G13_5,G13_6,G13_7,G13_8};
                                 sub_size*13-width: g<={G14_1,G14_2,G14_3,G14_4,G14_5,G14_6,G14_7,G14_8};
                                 sub_size*14-width: g<={G15_1,G15_2,G15_3,G15_4,G15_5,G15_6,G15_7,G15_8};
                                 sub_size*15-width: g<={G16_1,G16_2,G16_3,G16_4,G16_5,G16_6,G16_7,G16_8};
                                 sub_size*16-width: g<={G17_1,G17_2,G17_3,G17_4,G17_5,G17_6,G17_7,G17_8};
                                 sub_size*17-width: g<={G18_1,G18_2,G18_3,G18_4,G18_5,G18_6,G18_7,G18_8};
                                 sub_size*18-width: g<={G19_1,G19_2,G19_3,G19_4,G19_5,G19_6,G19_7,G19_8};
                                 sub_size*19-width: g<={G20_1,G20_2,G20_3,G20_4,G20_5,G20_6,G20_7,G20_8};
                                 sub_size*20-width: g<={G21_1,G21_2,G21_3,G21_4,G21_5,G21_6,G21_7,G21_8};
                                 sub_size*21-width: g<={G22_1,G22_2,G22_3,G22_4,G22_5,G22_6,G22_7,G22_8};
                                 sub_size*22-width: g<={G23_1,G23_2,G23_3,G23_4,G23_5,G23_6,G23_7,G23_8};
                                 sub_size*23-width: g<={G24_1,G24_2,G24_3,G24_4,G24_5,G24_6,G24_7,G24_8};
                                 sub_size*24-width: g<={G25_1,G25_2,G25_3,G25_4,G25_5,G25_6,G25_7,G25_8};
                                 sub_size*25-width: g<={G26_1,G26_2,G26_3,G26_4,G26_5,G26_6,G26_7,G26_8};
                                 sub_size*26-width: g<={G27_1,G27_2,G27_3,G27_4,G27_5,G27_6,G27_7,G27_8};
                                 sub_size*27-width: g<={G28_1,G28_2,G28_3,G28_4,G28_5,G28_6,G28_7,G28_8};
                                 sub_size*28-width: g<={G29_1,G29_2,G29_3,G29_4,G29_5,G29_6,G29_7,G29_8};
                                 sub_size*29-width: g<={G30_1,G30_2,G30_3,G30_4,G30_5,G30_6,G30_7,G30_8};
                                 sub_size*30-width: g<={G31_1,G31_2,G31_3,G31_4,G31_5,G31_6,G31_7,G31_8};
                                 sub_size*31-width: g<={G32_1,G32_2,G32_3,G32_4,G32_5,G32_6,G32_7,G32_8};
                                 sub_size*32-width: g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                                 default : g<={{g[sub_size*7+width-1:sub_size*7],g[sub_size*8-1:sub_size*7+width]},
                                               {g[sub_size*6+width-1:sub_size*6],g[sub_size*7-1:sub_size*6+width]},
                                               {g[sub_size*5+width-1:sub_size*5],g[sub_size*6-1:sub_size*5+width]},
                                               {g[sub_size*4+width-1:sub_size*4],g[sub_size*5-1:sub_size*4+width]},
                                               {g[sub_size*3+width-1:sub_size*3],g[sub_size*4-1:sub_size*3+width]},
                                               {g[sub_size*2+width-1:sub_size*2],g[sub_size*3-1:sub_size*2+width]},
                                               {g[sub_size*1+width-1:sub_size*1],g[sub_size*2-1:sub_size*1+width]},
                                               {g[sub_size*0+width-1:sub_size*0],g[sub_size*1-1:sub_size*0+width]}
                                              };
                               endcase
                             end
                           else /*后级模块不能接受数据,本次信息位输出未被后级模块取走*/
                             begin
                               s_axis_tready<=0;
                               state<=STATE_waiting_ready;
                               if(s_axis_tready&&s_axis_tvalid) /*本次输出未被取走,即使输入端具备有效数据,也不能将其更新至输出,只能寄存*/
                                 begin
                                   s_tdata_reg<=s_axis_tdata;
                                   reg_flag<=1;
                                 end
                             end
                         end
      
        STATE_waiting_ready : begin
                                if(m_axis_tready&&m_axis_tvalid)
                                  begin
                                    check<=check^check_reg;
                                    if(in_out_cnt==k-width)
                                      begin
                                        in_out_cnt<=0;
                                        m_axis_tdata<=m_axis_tdata;
                                        m_axis_tvalid<=0;
                                        state<=STATE_check_out;
                                      end
                                    else
                                      begin
                                        in_out_cnt<=in_out_cnt+width;
                                        s_axis_tready<=1;
                                        if(reg_flag==0)
                                          begin
                                            m_axis_tdata<=m_axis_tdata;
                                            m_axis_tvalid<=0;
                                            state<=STATE_waiting_valid;
                                          end
                                        else
                                          begin
                                            reg_flag<=0;
                                            m_axis_tdata<=s_tdata_reg;
                                            m_axis_tvalid<=1;
                                            state<=STATE_data_out;
                                          end
                                      end
                                    case(in_out_cnt)
                                      sub_size*1-width : g<={G2_1,G2_2,G2_3,G2_4,G2_5,G2_6,G2_7,G2_8};
                                      sub_size*2-width : g<={G3_1,G3_2,G3_3,G3_4,G3_5,G3_6,G3_7,G3_8};
                                      sub_size*3-width : g<={G4_1,G4_2,G4_3,G4_4,G4_5,G4_6,G4_7,G4_8};
                                      sub_size*4-width : g<={G5_1,G5_2,G5_3,G5_4,G5_5,G5_6,G5_7,G5_8};
                                      sub_size*5-width : g<={G6_1,G6_2,G6_3,G6_4,G6_5,G6_6,G6_7,G6_8};
                                      sub_size*6-width : g<={G7_1,G7_2,G7_3,G7_4,G7_5,G7_6,G7_7,G7_8};
                                      sub_size*7-width : g<={G8_1,G8_2,G8_3,G8_4,G8_5,G8_6,G8_7,G8_8};
                                      sub_size*8-width : g<={G9_1,G9_2,G9_3,G9_4,G9_5,G9_6,G9_7,G9_8};
                                      sub_size*9-width : g<={G10_1,G10_2,G10_3,G10_4,G10_5,G10_6,G10_7,G10_8};
                                      sub_size*10-width: g<={G11_1,G11_2,G11_3,G11_4,G11_5,G11_6,G11_7,G11_8};
                                      sub_size*11-width: g<={G12_1,G12_2,G12_3,G12_4,G12_5,G12_6,G12_7,G12_8};
                                      sub_size*12-width: g<={G13_1,G13_2,G13_3,G13_4,G13_5,G13_6,G13_7,G13_8};
                                      sub_size*13-width: g<={G14_1,G14_2,G14_3,G14_4,G14_5,G14_6,G14_7,G14_8};
                                      sub_size*14-width: g<={G15_1,G15_2,G15_3,G15_4,G15_5,G15_6,G15_7,G15_8};
                                      sub_size*15-width: g<={G16_1,G16_2,G16_3,G16_4,G16_5,G16_6,G16_7,G16_8};
                                      sub_size*16-width: g<={G17_1,G17_2,G17_3,G17_4,G17_5,G17_6,G17_7,G17_8};
                                      sub_size*17-width: g<={G18_1,G18_2,G18_3,G18_4,G18_5,G18_6,G18_7,G18_8};
                                      sub_size*18-width: g<={G19_1,G19_2,G19_3,G19_4,G19_5,G19_6,G19_7,G19_8};
                                      sub_size*19-width: g<={G20_1,G20_2,G20_3,G20_4,G20_5,G20_6,G20_7,G20_8};
                                      sub_size*20-width: g<={G21_1,G21_2,G21_3,G21_4,G21_5,G21_6,G21_7,G21_8};
                                      sub_size*21-width: g<={G22_1,G22_2,G22_3,G22_4,G22_5,G22_6,G22_7,G22_8};
                                      sub_size*22-width: g<={G23_1,G23_2,G23_3,G23_4,G23_5,G23_6,G23_7,G23_8};
                                      sub_size*23-width: g<={G24_1,G24_2,G24_3,G24_4,G24_5,G24_6,G24_7,G24_8};
                                      sub_size*24-width: g<={G25_1,G25_2,G25_3,G25_4,G25_5,G25_6,G25_7,G25_8};
                                      sub_size*25-width: g<={G26_1,G26_2,G26_3,G26_4,G26_5,G26_6,G26_7,G26_8};
                                      sub_size*26-width: g<={G27_1,G27_2,G27_3,G27_4,G27_5,G27_6,G27_7,G27_8};
                                      sub_size*27-width: g<={G28_1,G28_2,G28_3,G28_4,G28_5,G28_6,G28_7,G28_8};
                                      sub_size*28-width: g<={G29_1,G29_2,G29_3,G29_4,G29_5,G29_6,G29_7,G29_8};
                                      sub_size*29-width: g<={G30_1,G30_2,G30_3,G30_4,G30_5,G30_6,G30_7,G30_8};
                                      sub_size*30-width: g<={G31_1,G31_2,G31_3,G31_4,G31_5,G31_6,G31_7,G31_8};
                                      sub_size*31-width: g<={G32_1,G32_2,G32_3,G32_4,G32_5,G32_6,G32_7,G32_8};
                                      sub_size*32-width: g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                                      default : g<={{g[sub_size*7+width-1:sub_size*7],g[sub_size*8-1:sub_size*7+width]},
                                                    {g[sub_size*6+width-1:sub_size*6],g[sub_size*7-1:sub_size*6+width]},
                                                    {g[sub_size*5+width-1:sub_size*5],g[sub_size*6-1:sub_size*5+width]},
                                                    {g[sub_size*4+width-1:sub_size*4],g[sub_size*5-1:sub_size*4+width]},
                                                    {g[sub_size*3+width-1:sub_size*3],g[sub_size*4-1:sub_size*3+width]},
                                                    {g[sub_size*2+width-1:sub_size*2],g[sub_size*3-1:sub_size*2+width]},
                                                    {g[sub_size*1+width-1:sub_size*1],g[sub_size*2-1:sub_size*1+width]},
                                                    {g[sub_size*0+width-1:sub_size*0],g[sub_size*1-1:sub_size*0+width]}
                                                   };
                                    endcase
                                  end
                              end

        STATE_check_out : begin
                            if(!m_axis_tvalid)
                              begin
                                in_out_cnt<=0;
                                m_axis_tdata<=check[n-k-1:n-k-width];
                                m_axis_tvalid<=1;
                              end
                            else if(m_axis_tready&&m_axis_tvalid)
                              begin
                                if(in_out_cnt==n-k-width)
                                  begin
                                    in_out_cnt<=0;
                                    check<=0;
                                    s_axis_tready<=1;
                                    m_axis_tlast<=0;
                                    if(reg_flag)
                                      begin
                                        m_axis_tdata<=s_tdata_reg;
                                        reg_flag<=0;
                                        state<=STATE_data_out;
                                      end
                                    else
                                      begin
                                        m_axis_tdata<=m_axis_tdata;
                                        m_axis_tvalid<=0;
                                        state<=STATE_waiting_valid;
                                      end
                                  end
                                else if(in_out_cnt==n-k-2*width)
                                  begin
                                    in_out_cnt<=in_out_cnt+width;
                                    m_axis_tdata<=check[(n-k-1-in_out_cnt-width*2+1) +: width];
                                    m_axis_tlast<=1;
                                  end
                                else
                                  begin
                                    in_out_cnt<=in_out_cnt+width;
                                    m_axis_tdata<=check[(n-k-1-in_out_cnt-width*2+1) +: width];
                                  end
                              end
                          end
                          
        default : begin
                    in_out_cnt<=0;
                    g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                    check<=0;
                    s_axis_tready<=0;
                    m_axis_tdata<=0;
                    m_axis_tvalid<=0;
                    m_axis_tlast<=0;
                    state<=STATE_waiting_valid;            
                  end
      endcase
    end
end
/***********************************************************************************************************/

endmodule