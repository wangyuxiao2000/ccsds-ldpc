/*************************************************************/
//function: CCSDS-(24576,16384)LDPC编码器
//Author  : WangYuxiao
//Email   : wyxee2000@163.com
//Data    : 2024.1.24
//Version : V 1.0
/*************************************************************/
`timescale 1 ns / 1 ps

module encoder_24576_16384 (clk,rst_n,s_axis_tdata,s_axis_tvalid,s_axis_tready,m_axis_tdata,m_axis_tvalid,m_axis_tlast,m_axis_tready);
/************************************************生成矩阵设置************************************************/
parameter width = 8; /*支持1、2、4、8、16、32、64*/
localparam n = 24576;
localparam k = 16384;
localparam sub_size = 1024;
localparam G1_1 = 1024'h2A1944B6A513DA9A23E91B538352D9051D55C7968FD8B60DB12C8D35E8B947C57FDAC5E20E8E406043C56EF199A6CC68FBA3C2753FAE011BDA4E5C55F45164C187292033229B6AC622263EFE363002769C0AC7E3735F6D6A6064B23588F9C7B22311DB8B7A0015AB60998B1226AEC289AD36CA4D9A0B4E147D21C1491E9F601F;
localparam G1_2 = 1024'h582FA8B195AC0FF6B17494C80D7D3103538D5CD4158D7016EDE15E90A8B991A7E65531FC88C80C53F50757E3C1DBA4A9941CB9E10CA85D4CFAF32ED70F835F5C34957AACB36793F1A60D8D589ED970A3B709D10A26F0AFB4278635F21C5E303BEB168E59A4F8186B2365928C6EE6C2288944BE90042283A84237F5DACCB99911;
localparam G1_3 = 1024'hC402CF86161B7FD658999EAE801FE784ABFFF14E49D1DE40E531BF3B0054BB38C2C19BD09D2DC2A0565B95CE5B09AC3659E7F519F7E0AFA778EE264848BFAC1873DE56D6916CD06E1517435E10326FE1FAF7E3A5B9E94FCF64390AF7C713374DE1CE8B53AF3ED21F4491D46179014FC0B1CB6A4877FD296000B1CD22B137AF9E;
localparam G1_4 = 1024'hEF7FF4F5C55C2176A91817D8C1C96970A512A6EAFFD60E46109F98FE464AAE2747B9DA6031E5B50748B9A2EA8E88887A138E243B8D213ED44DDAB36219750BE09C4C54F7AA8C7F12217CF431E0D23AF414817E58ACBCFBF8C08ACF0D81D764ED395771F769430700C6AC60DE506F75820EC751DE8FB8056841B6B7A2540C5EAD;
localparam G1_5 = 1024'hA7FB9B612C519149BD93961EDC8759F3B8099F669D56F87330F65157087A86E44FDB481C90599168CB3E93B5A2E4511D92E2EE2BC4CA1E64F9D040608C5AB3B75C9F7B484797F5FA389577CDE7FCFD8D4CF0C5FF7848297FAFCD479F55382A4D6F965B93B98AE8710E3D145F20A66698AAC31BE86915568980F8873EFF01AF6F;
localparam G1_6 = 1024'h7A9675133B748526243F7E24BFB12FF0F00FE99253C417C0598B635414E65035C84D6C17CEF34D71CDA491F3A4CC61311CAB65D743C7525D25FE6D8EF17C5EA64EBD7558B5B37B54E6CD260D58FCCA11E495DD026C0D1750F3083AA6C785DF66975F4E955111793A8713F0A7DA83FD74260D7B929FCC46247F5BB0A475B7328F;
localparam G1_7 = 1024'h7B927E11105C995F4C95736351CB287B0F27D794E840EAB57CD1742148459596A533EEE84463C707B418F663B936EE7C4F73B1B2EB99E9216FAA2F137DE9085D9C097D3F33128DC844ED946F943DED2EBFEF4B7B1FD1A721D13A3691A640B9EEEF40A4B21BF9D397A3281F112B4BA26600FF74F713124CE0EDED3B7DE98C35F4;
localparam G1_8 = 1024'hAF11E6E8CE5EE091C8E64FD90B593DD98003981EADB08B189F3EB25FFA593C49D76C1A21B1DE760196F9375B617E3E8CF5729C7D1656BF44EB5003F265B89151DB13557986503EFB28448ACDED78EB00E40518751F8330A20409789A67390A87D72CF3BFEF98B57E475628890132F0C29A7CA2BB3184BC35D8A963010CFF7C9E;
localparam G2_1 = 1024'h849B64C14825CA366FCB6F9B74AF982AA35F4CA37919A32A83988B6A6623F245CAA4043983F2D08B3B18BED0284154D8BB3969DE8D3C668F5F0FEB22536F42B0D6AC347474B14CCC4E87E418327EBBFDF0618019610390EAD3D53291E457D2D3015EA4900D216C19969E52D88FA512712CF7502FA4B95F230226BEA7DEE79C0C;
localparam G2_2 = 1024'hB7E065CFEE395036DF10295F9B2C93DFC5F718ED209ADCE32998A7B3B8C14654C1341FD42A2E9A710D7BF1717BA9D0E6EB69F20722BC59ED79CF45BA8C3C47F4BBEBF615B6BDC20483B47A96C9D34664ED8513E9095A74E2A918110EC231E26C8695BC53AAD7F7EDDF9F9F6D228AC2BEB4FCC48882AD371C9640F612C559DA7F;
localparam G2_3 = 1024'h00F85B84D77B53ED8E8BED5D6AE55252CF92A4B1A5C9A979B3BBD5CC2BE97C2443AA2DF6B5252F5967C1FB678EA8163FB86DEA872FB8AD09551F3C7FF3FF7FB2DC1F38F020EE532EBFD791636110D31D1ED811C5E5250AD86255C718F555200619FFA9C1565EFA23B17D8C1226830A763CC442A9A5DDC77E4EEF6FB39F069B41;
localparam G2_4 = 1024'h904B9F993776FB3041C8AD9B1618EFD4C31840CBB79B2F5FE280E48EA3163A5B07809FDDC12D6DB186A59371F1586F2F7B4D3F67FB7B90CBEC97C751690E0C666D647DED3F065BF571552047A1736C0CF2C68E0D898B924742863937C0BB2611BB7771237B3B44316881CE1723F58ACA7E4F423D03C31394CED6FBDA27408A61;
localparam G2_5 = 1024'hCBE42896973658B8BED649F09E51833935D9DE3AF89FEF13EA78B56806964505BAF2922A27587D56D1DD119C138FE30FD7BA9B4F9FB638DBA120449568571F6B483A2BC9FC0BA5685C2FE1E9BFE650E6FFFAB3498592BD3329AC0C5E4AC0AAE54634A1F964A8B5DC243CA901FC281A13BEE0BFB975F01D37335A442227E3EB0F;
localparam G2_6 = 1024'hECA9294F817237DAED7133CAF7245C3269A4E1CFD6D553579579033C94907C6F3C24090292F165E1425F784FC2E4DC130BFC4155DCAD777AB3E54CCE726B7A9D5A99EA132096D34DD4AE25E971B834A4435E940089B047DA62A9D11D3F7997C927FFFC6F61CDC4342C0814DBAD8BE04A9EBB8A126FD6FEFE5602B1B5A9A2E355;
localparam G2_7 = 1024'hD810242CC8CEEC9B2A435E01970CEFF4D92C23C480C827B285F81BFDD54C0853FE10BD450A5B52EDEECD89FB768D8DA0A9BE8DE517A695B16CEAC36C8638E1279EFC71D26B7D11D50577A7E6E586D098400D7574D4A696558D3DB1A8D9D843C788C7694952104975647D6DFA3DCEFB416E6AC77F562AFA47D30A1DD983FB332E;
localparam G2_8 = 1024'h3B55AFAEEB396DFE102CB12B0C22B21CC11AA85369302814AC4A5E85E020001FF902E721DDCC5DF9D9AA63C438E0C3AE5223173A822506689C6C71772C6D9AE6DFF95978C6552A1A4E86AEA19A16249F9BE1ECD7AEECC01CC3BF4852FC784342B4A93D0B363E81312E893951B8E4BA431B6469A8E686F962CD39F0F590F0CF76;
localparam G3_1 = 1024'hF1EF407C6F6F4233133BD4815CFB10E96544F957495D52BB9654321C2ECC9883A990726F052D8ACCC37DC53FDCB5E2B4FE2E70E242CCDDC5AB37DD64E9087014836ADB986B84ED3A078101C832BBE0097928F249CC69EA20A02C9AC575386B7CFC0CE60B8BFED1381057591AD420A5543EB1C3D419CDC5A672F25EBE6EDEB835;
localparam G3_2 = 1024'h889A6B1934F029DCA63C61DF31DEF89DE1911403BC0BF0B53D0DABC81EC3C13CD048A302D3AA739E666BA3A62A2BD58068B08D0DB9DF4EB6512407995C00D194986384BBDC575FE580FCEF34E1E25B606E8FFF39CB1399F655B36CE61EF37C2F50C4F3732283482DBAF67B1C7B229D677E0409D0D7762F17C6DE4F97C402CED5;
localparam G3_3 = 1024'h7751FFD538000D8BB70D7C48C459E3B816F0E14C9572067575C64C764366B79471C95F606C99447E6CB89458D1810951FA11CDC92BD810C4D41688DE35C17602D3229C338D4B2C6D9D8A25C88CAE544C968235191802D83ECD088AF24CD2BFE877092C5608C335648737CAEA1E0055CA80897A26C3A3615119AE8D8A9D6EC8BD;
localparam G3_4 = 1024'h384802615179A68E94C16A7A5B914847CED75D4C913F0055102C49E0E1636371AC9A6298928FF649394C30C59EEBFF5EA8525C13D9A1FC21629D2CCC80792CF66B482C7E6E59599A9B7854E6C2492A29F5047C8075A8F1218A8D5BE016636D61860D274C0EF3749EADF2902F09D221C534720ED4F0DEC03020DCF5BF3B8640D1;
localparam G3_5 = 1024'hA815CD0110EDAB82DDEB86277E006E8947632CACF7C15569E98E167C38F670A1E938F6E64A75D4F0F0647E493D27845FCCD4CE75D0FEBE8C7CE78C25EBC00E54A6592D4C375D1475E1B331922024B49B82112F4F4CF7966595AF45FFB1DFF7D7AF283C8C75E2B4EBAD82D4C002F678BC2FA8206DF324B10DA06A635321D1897F;
localparam G3_6 = 1024'hB8BE6D489F5ECA6BF0F8A470BDF10F0E6910EBE3D47D63FED1B1AD1411ACF684943B96E33F14DD2CCA7A18120F329616CF2DE7E47BB21A122F688AE2404FB6DE449931DE1B7D1F435CB5CF80F591644FF891BED8E3DA85C3DCA903F2D75E3E2DC7DF7DB3EECBC2AF485958C608150ECFF47B6D612827794451C8CE43604FE3EB;
localparam G3_7 = 1024'h338A85E48C3BA52DC6EC976BF87F68953A5F7BAF0482FC7CBC487E99F0BC51930B11116A9A8EB28A02F7CDE4300747EBF995466FB729E7FF0DA2C3CB00258303353765881788F8D2D777C56973BB8CCE28CCA2161D3785BE9D62839E8702A4BBB125FBA16BDFD2689100C4084CF678DE28442E1159562F42A5753C53B02C4395;
localparam G3_8 = 1024'h56966F31B8F46D9598B33E134BA37F5E8D2163A0F33A1EA1A1BB7E0776DA6D05AF5B92172DB479D82C2B23868D90F8F6000D8ECA22EEF0556C6D11B8803561FC508DDFD60520DC939751DC3BF042FB4673BAA7548275279599297F4C96FCF0039A419386D4E73749DA479DBE3F7BF61537F3A9487BCFB090D159370A87911D17;
localparam G4_1 = 1024'h5F418FC3CFAC0C53F665AF0AB3DA14725DDE7F677681713C6C8FCD921D6BB5FD3AF9FF06B8F070759AF26FE23CE6B984D8227A4EFA4673252B44A6B59AB980C7E4490288B1A148C7D5B1093B080E43BD0B36828C33C6215B8DB290D6242B0A0AEFCD377EA2DDE7C401D4CA015900D13C797C702E2364E2FC9F90C19D36AFE361;
localparam G4_2 = 1024'h7D4DEE216BAB3D95CA20D51EDF295530B16A08192A7AC96012440DB6BC5B530C86F5CD8BF6023CAE582098AB7FD61E9AC10919BB205D25C105A44F798748CC4230EA5AA24209DF6016E713B3AD7908BC89BC44F15132762DC37E95A0E2F9EA38ED60FB2368C65F3E4439BEFA80D80276EEDEA0A8A64911000DA4D5B243908903;
localparam G4_3 = 1024'h316181AC4642C974CFBDFA8EC441F921C1EB801CA85A096A572F605F2B27DD559A1239999C1263BA3D119ABEC0E2CF9449649686058BE3752FA129FEBC88FF17218292376FEA74ADF23FD0DC7D3E66038F618DAC28F4D4070D8B02A6BE1ABF9078E672B4C33BEB2B15A7DD62670A61BE4432D7CF2F015C149F133D901F9BD2BA;
localparam G4_4 = 1024'hF3A8315B315AF888C0C399610BEA4CF019C830BDD0B08D0A872B01547A5280FE83F4F8849C09791425282042B408428F7705338DD026798DE5997650C1331A9AD9A4A7CB073D4C32AC2C5737FE15F0BE3394769416B1FFBAF64B64FF364544E07DBAF47E432CAFCD7FCA2B48F0432466212F6310C4782BBB759E894F5D7A498A;
localparam G4_5 = 1024'hB90806CFE206D9C8C667680CC9DD4BAB94B3A49C2F7FD82743FB1F22AE4BDD7C43F9868D6802192369AD5377762593676AC81BEA3F3AD0003572B7F3C39BEF8145193626BB96378DAB46D3AA32E8CF14CC0400337F583D4C090A6204EA76B9C88847F648163AFFE20B8F2F100663EF61A8EF2C23EA933B41DA49EB24AB53A9A8;
localparam G4_6 = 1024'h5E96FBE090B1282D7D77B46C962C0087BD4C4F5E5C583AEA90DD7BE3E531B27BC9A6FABA0A32668829C56A807C1012DC2453F15A2A1ADAD904A9C5B0CFBF4C36B845C3D97FB5B5E0495490B897B3FB90EF4D318420297BFC027363DC92690F76478C4E0752E03BE3D2E86CB59084124C1E6C6A3C8A159D1ADB0899952915E695;
localparam G4_7 = 1024'h731399C402086762EBD25F0DCC505D8EEA7E44CAB4D351C0BDC7FB3A12EEFC9F26CDBA52F0A011607183806E4F8188B205D3D58A46D21B6A4A6AFB84015AE156FF63A4DB65D6975CF70B62C40BB97C887D7584DB8B4EF722DCA95C7D070A1F4F197381F7848E80DD2A78105BAE4B512B240CFB9F147BF27399142CB9E5FF2BF6;
localparam G4_8 = 1024'h3BF8A96B457D6B93EE72DECFAD451230C4D30C7A831824B494D8079BC28B93534C37DECA1DECE16237F4C4555AA14F7FFBE8733C2FCCCDF75432D88765504FA64FE2E4F9E410765C4F8988E12889B368B97B2D9FE9E56C35410C9959FCDB43C05E45882F985798F7331A76E720F29295D6AE7ED0B26182F7333232901582D1DA;
localparam G5_1 = 1024'h10408E1CDEE38759D68341099699860E6361B870B4C461274229F0B721D0E971F1027AB653BCD35AA72F6284780BE3322F6AF953D13F6ADE5520F200335FA0C24DC6A54DF45EE2A6EC1FBD0EA5825AF4AA7AE4473EA69EAD8DDB064E9DE08E5E8C49B32D75726282E5745021728D4F868253896F03518263BFDBB6A0FB6A9485;
localparam G5_2 = 1024'h99C79A8CA490E24CFC2B61BD417C25F76F4C435122526720F52774D99310E74E86F74AB07231D7159FABF13B9383CBD9D45A7E375AB534774250E4E8452D37623E651AD302A4325800CD7480CC10AFD1F9AC7C628587F5D6AAE3C010866E42E85E9325176764B4B1B52C6C2EF2021208D4260999A207967FD43B77788D37FDF9;
localparam G5_3 = 1024'hACC128EFC68E2A0B73477E1B8F3536A10D578B55FEC4C12031937B1C73D05640B93FEA661F10E57886A0407E643ECF561AF56B703AF0F24314A332F8F5ABC11881ED24B90E9A0BE991BEE2E4223A0B05469CA8CB6AB1DF0C805C6395A995DDE44380F5FFDF9373B68BFBD1B3B3E7C7E6291D20F32658F56D29FDA8C44EAC5EEA;
localparam G5_4 = 1024'h193FC68594530A894C0F9E40F23F624F6E60D786AF2466845CBE5A553F574416268AEF9F12689E5708093EB40BF289ACDD18AFB31CF2217508F680F95748112D5A94EEA3D8940D68C7418BB34D15AFC3ECF0A71BE0CC4F42B719E5ED9E0F4DF279426319DD0322E1C6421792FC8E51A951B0BB5A7EEAEC214E8CD4E5C12DD232;
localparam G5_5 = 1024'hB40B27AA43F555385A0B14438FCA941E1BF19878880DD1D7DFCBA051C1BD370447B7BF271F2B1D07DC6687C1764B352062BA1957EBBC1A19214F49C843F701086DE3E22963F7E0F1888118670EA15BAF3BE590C9CD1BE8A9641E43D842A7D2E9986D9D74512593147D7FD74D99B736861656AB9904B648B39121932A4CFB809E;
localparam G5_6 = 1024'h5B59F58D4AA4BEC2A1A1FEA7D7A0A6BC04527680A7F6456AE41DBEF103E456FBD2242146AE879AA50C04F67B92190E80139FEA972A1A21EAE45A88298E32FABB4F564FB195CDEF4BB0CFDECA8BBA1139ABE26DD394F0A68806A5CE7F68175B7D7CA6789DDE52A59DA4E64613DC81442F25AE0B6EB16355858D4F9A916A079365;
localparam G5_7 = 1024'h0306A55B4B9B4021C50EB6DC48E0695C67D1078F88EBEF99D321D1F7FBEAFD8A7D633DC23965273DD7C9587B27C29D3B428600ECCF1A93387E41DCF3ABD7325104437EDE0A8E465DF6EF9E247FE59A492B649919838693F8167A7572D5E34EAC5425D24622BB3204371A77A6A5E34BB4FD365D2F016CAA9938414F8CC35C1C10;
localparam G5_8 = 1024'h865C262BFF92F81C5588F1F4A53DFA4B3B8C3EF085CB59963E18E6AF366A0C07A0204795BBDCA4835A356A95BEEA8D21E53EDFF37D77A5CC3D051C6A0D07D6E5749B5B2FBDDCC600744A1981FDB3BFC3E58EEA88B6803F6FA66321A2620E8CEB342D02DBC212A28FEE9CECC1011699E71882D83851A3D97D647866242B9BFC1C;
localparam G6_1 = 1024'hB3C024A6D45738BE15105F83DAFE2292691E004B047E35B06C0353280BB1BE07D17E9BFF9A4879783C080C6875976CED517ADADF4CA0C4CB863938CC99B94B956F4DD9BE0161EA789F9AC215F2D19A3EC253015EA3FECAB7502089AB2186760717F558F73B58053E3B5E7872E772336B05D3977FE664CD172F9AA5E1373BB533;
localparam G6_2 = 1024'h6EF819CC4FB0F231401AD371DB38587FF1AD36FAD52985CDEB07FF0BE58540B093EB3319B9698EC7AC6C1F68929DD80C79173DD6F373A7439CDC071D84BDFE5B96852FEC83D971EDE842FE39470025514C47B9E3E1FA6690838484B3AE38883145FFD41A8347067C73E0D514D1430AB1DBC92D309325CD29BFBD320B75296C32;
localparam G6_3 = 1024'h6DBA2F587863BF99F4FA9B936B692E0FC14528780BDE33E318F290E16625CCB511472B57D5D27B5EE737A6BDCD5D7D130D56BA323D31A88F16B9D8829B97BAE254F5C49CAD7DEBEBE75800963C123757CC4AA38812D2CE8F9529B1610453549A9134679DC25459261294EBF00516C21BDBBEB30C0F86FCCF1DA682C21D9F6642;
localparam G6_4 = 1024'hF0E48C0A2021C9F5D86D16FF89298964CD0B301905DA47238935BA3F63067601F7A58F3AE5297F1BD628ABF7C893762360F81FC3803BBF077D7A20F8425AD62BE65CDE27CE457DA0EF9B239314F0B0BF1F5CC2F1169F45A50B971DDE2854E11B640D7675EE18A8ABE29E78A01CF2FFDA0E6937DBC60BBE6B40F08038E757B59B;
localparam G6_5 = 1024'hB3AA688B7FD431EF8D77271FD227AEA1F6534CDCDBA0CEE0C6A673F43986EB96C4CCC76FA65E02CA3419A1CBC02E3448125E40D5C455610E84196D665370464EB78EEA28DE582A4597A2DA98CDBEB1A2C77D35EFE90AF8C3FC1769F4EFF89931AA08B69BAEF31564137DF4737B24791BFDD583D5523901B85CE2E4D07D2DF46F;
localparam G6_6 = 1024'h843BF69DE565A4A7A8B716620C9815838C26E4B83B9435B76C38B28E0DAC28F124E4158A2F4EEC9D067B3A071BB48AC6D49945FBF1254160DAF1BEC7017843002E3F4D06F76CAD0CAAACF1041348471BAB17F5316B95292B01CB8FABE99062D4BC9968A8437E371AEFCDEEFA7DFF3B809587D6AF8F87569C015CD05ECBA23D8F;
localparam G6_7 = 1024'h355AEFA00B91CE52E5FE7B3443DD0EB46F39C0623DAE7398612D7050886BBFF853639ABA847BB032122EFEC43D5982782CFCB8B518B6A7AFA055550D57A25CB3453E083E4CC6CFE95B3C6B83547049E3DB1A8B63C17BA5E3F26240E0D849F0CA019E67C22A2E70B8EAEF37D58FEA7C35BE4FE4FA6005CECC3643674B43C06D6A;
localparam G6_8 = 1024'h3D6B3ACDC6DA7F47F14A05DEF18DAF79D9D2E5FB39FEF16B73BC0100DFFEAE9BCA1AFF9CE441BDC275821EF00EBF85B0546362CF2F45B344A56820B449C864262DCF43BE4BE5E35FCCA1E38029CE34711AA16C20B12A0853248AD295147A8A44F66C46EB7320B231709D0AC7DE68224CF638B4D87DA46773D0DC0BC12D440101;
localparam G7_1 = 1024'hA8B9E1E450675AF58036340DF0FC2B8E6CC46FEF366830A6F9537C4841A9AE514AB4372F672F66CF72E52311EA0C74298C36BE8CDE824B9238ACA030934D005AB2C67BE070D15B3830E9AF3CD07A57323652EB1FAB2FBD786DADC3C2C467ED9E34325C805C6D7494C329C1806A36154949547DC04262E3E20103B93A0E5E4B88;
localparam G7_2 = 1024'hBAA7B2BE7EEA13439C1D695F26233684FE8AD7F9FE8FEE4A05369494C1BEE63495F4F421F748781D0EE5B926036F457466685DBA4EC5F3EB6F6A4B85A0EB94FC89E21201228056210DC2C2EAEF22B089CAC880CD907BF162A908594B535932B3D41AB0C582E6253E37253A9FCC6727E97CD1421DA318D90FB54B061F7B53AD2C;
localparam G7_3 = 1024'h81107A7CBE1D769BBF0E2664D5396DC52DCE1CD44E10B816E8783409DC6C5AF51B81A00F9BDA49E66474F08E32CC2B5ED8A3D389C72F9EA4B8ACAA9A78C594BF9F50666FFDE24AE3FCF2334C3F571E2F29AE8AAFE9CB2C349987134C14D48631D9F5FD824C9A8BE301D6B3AFF57C3E4E896BF2A57C016B9C0E5C3AAB03EFD0F9;
localparam G7_4 = 1024'h85D2686AE0D1BB45173695244935699AB522A9849303E8EC5AC3835EDA7AD68DF76BB7D31A26571F423F79EF01E5141F4DFF64AE417C30094E6B1DC6B9318BE1EF9520A64BDF761307E01F114004ADA7EC7D92AB34703AC8BC71221CFB984E72C6DE69F87535D3B7E8D46C6EF919FB14ED5067638B48F14BDD7EFF6EEB0E774B;
localparam G7_5 = 1024'h4A612448249EC967138B7CE7110CBA054EBCCDCC2BC3AB29F32330541043A4134301ECE943D0BE20851CA8AE5CBBC1E4473A390BAC5D4C7A5C55FAAA26299718998488E16C7EDBE24A3FE798889AA4E4DB3B10D6D4FD86250229A3D1B53703B0FD600A04B2FC45BA0B9B11443B823B073836F95CD5E2D3397A85DE4E05829DE0;
localparam G7_6 = 1024'h5BF1EAA5488597D72B8AC5B844FE18FF34A7AD93E0B7DCCEC2259A6D96810AB631DDACA6D5BDAADAB521D561CE4E62766F8924057F2121CB72373B9887798B8FF7FD29637A9E1690A1199E6D90E4B8D354002F8B1349759ED192C7D62711F4B618FCB84889ABBCA5927053E73746896A0727363A64EEE4758D6E46E72FE76ACA;
localparam G7_7 = 1024'h22963EBB23E0AB094A1D24EB920C29C3676D60DA7FF24A2C7480E75F7F02E8F5F4C3856FF0F5BDF99AA4050A61BEB59437C8F4DFE371F647AFAAD2486CBE008A3A01E907B9AC0E8F876027409C9E1A784BD9AAAE4EB56FDDA7D94A571722A8078E30BA7D28D66E78A1015E0864AEA4FF59CA6179B8184D88BADD1956B35E8DE5;
localparam G7_8 = 1024'h8D55A6523B81C174B6A25773D7033CCF8096F33F43FB242B8EFF2EF7A79C8E8F878E8DEC27475DB895CE5F9A8800DE259FC4076F9D52579DF3FF8CB1CFBD94BA18C8B2FF2692BDC9A65E5982E12E04F134B4C5C459327F4D540090F2DCDCF6F8A4D7B9044DECB7793F57C655ABEA48BB5A26BCF1709A8039C63C0DA0872C77AF;
localparam G8_1 = 1024'h0835CA7C32ADC04B48A273B0A9278CC4B4E05B666419EB18A891F0F1FE75A5EE5DB0303C94181EC15A480D624D518BEDC8CDA450CE9566C683CD287C072B1CCB667BD82F14342209F0156DB27F74A37DEEF3F235EE26B4B07A8F1B281E9325CB6E9FA21672808C76F03687392364CDE646294FB4B2098C51E10C7B4FA32C0ED5;
localparam G8_2 = 1024'h634E9D5639336A928EFB2B1B32F44E9E1060BD198E5952B5A074A52C8CB82CD7C936647C9D75967A0C3B4A3F9ACFA548FD71A471DBC3560BB00894F0EAF37724D70C2A4130F2002B974D9619806AC2B076FE2E7DF386BD07FBC520810A19FF455E377B89D6549ACF6DCCC8D6593EB6969581394F65D885978AC7A63AE3BD533C;
localparam G8_3 = 1024'hE0AA5F1D3498290A6F47317417AF1A6F515C508B025EAA7F5C8A6D6FAF173A8897A64EBD6B7BB758447C486791F5CDA4799A07A5DBF3580EA1F92DF16936D3A10B81734C73452A23193AC1B64DA2B50E27ABB4AD9D1E4A5B5CA076908771181CF8D9CD0B6F4E17E3422BE1A45135F7483190A6C7044E3EBBE206388F247471DF;
localparam G8_4 = 1024'h2ED4B04FF33DA75A74C296D5236F12ADB2F9EF5BC8EECEE71A069E994E9EDB545759ABFBEEFC49BA3182A827C232E3518E9C30CC96ED4FD7232CB7C466E267C6343EA7069707D6D82EB4BEAED6CCDBC8402B41E6E25BFCF11E8CFBFCF26C749B7096D7CE94776FCC2FE3D084D6D95EA903BD4C8B6A57DFFA659B085CD1A298A9;
localparam G8_5 = 1024'h269E0458427E616DE7382E7B4F4F2FBEDA8BF281662F2E51E8794FF15A9901DB38289BABA63CBC489F67E121FA8730464FE0585DC3590D2488A60C84D37D5414C04519CF7FCCE12C34C0F1CDDC3DC5C32B36C6430CE624D6940F5239B3830D320C7C4F64B58AC9BEE203B9A6E9A5B5AD4E26B7ADFF09F2DF89CF907FB7A21305;
localparam G8_6 = 1024'hDF1F56A75C0FC4F8BEFE6A8A05E37CFCC1E35474745F2D00A781E922F543EC56552492C5D12F22311C6160144307BB91D11EEDDFFF47CF1ED79E2DBBC449C8C477515970CD8A38C7905762D4F22CECC610F087724D5AA56DAFE7595A62B61DDCDB2DC4CECFB548A6E20E11F6CDCB08D0CBC219EE522F246AC43BD8867061352D;
localparam G8_7 = 1024'h7ADD886B26827B0246240277B694881FAE72767976842858C0FEDCB1F7238B790B74AF64BC1D56C54089D5AAB6A71CA64F7E0DE8618CC14FDD4198F04C9DCB98E3DA8A79E0DBDFFCEC33D9ADBB934303C658A576A9C9D086D31A6E78A0B3AEC8576FE459E8023770716F38EC8AC4D9444C690B6CFD7428957E35DDBCE8524285;
localparam G8_8 = 1024'h59B63A6DD6940758B1C75EAC81C3EC4A284C88057A67ED8A6FACB5E440781D2DA864091B8165433C49C039F4FED29DCCF4BE8051FCCC3DC4CB4B56383DC6A052649A46BA038D2DAE5630DD5D178DFD00770E9F43197B22575A0A286009719192E0E9515708ADD9FF0A475DADCD586A007478D43F57996147516942935499F9BC;
localparam G9_1 = 1024'h0E0391250DED03B3CD57CEC1978728602020BB8AAA98096F53FB2DF7A9B7F76EC4237B1CE72541F26DBBAD8238E7EA4D11DF7F3F9228B8FD190E9EE6ADABEED176B7F2D56690DCD439D5B131C73A1714ABF442783A8DDBF0294215C58BFA0938AF9CE1D989330C518E32FF60C1517DD0993D6C233C3B71509C3020B95C2CA7EC;
localparam G9_2 = 1024'hE2072B04AF078EA5F49D3F6C2576C38C0740A72546C2BB02EEA51AC4D58736D5B8AFAC76214C26DF71FCD5A76E5AB65B7901D32BB89794478088E2C887F416A3CDC6F983E8444067A9E37129EA547EF5043ABDE86F20ABFCDCE105BA77DEE426AD8DC9FDD9A266E8FFF79B3F69C20CD76F893A0025C9001EE8D4550217715D82;
localparam G9_3 = 1024'h57D5322884BB4B7CDF7616A5159AAA641704AEE99603114B8CDA8BBC97F6E24005CB47F61BC076B5DB6345A333696F680E9D9654098DC12C7517D62267F6CB26AE9BB361757C3513FCCCD5E030C6F547E15A2EFD4636005B2CB33D9333980F11CE46E6E1568EEFA7B0C3A73EECAE13229D78435D928E00F62C340C46F25BFA19;
localparam G9_4 = 1024'h7C809C416C9D6A9BFAECF1DB2B4B7CEB4C5E98DA074FD752E322C24FD1258F9003396903A4C5AC59FD8B67AFD3007B0CC4301DB850BF6C6F9EBFF01CA092B7A014531DA7A1C5510FA9943875DB1855291B0AFD3A2359B545E90CC68A3FEC07E7D9199E2E8DBF3AF6141AF66A3DC869FA2280D00DEC92F9ECA768EDEBE61621CC;
localparam G9_5 = 1024'hBA34D42DB9A5571FCB7033BEF7A04128182E74BE31907455A2B866DB33A1982A9805B7C5CCA7F8E4275AB956264D2258C0712B3320837DEAB4A2F75498EF05FBB729B958B855D4606C6648EF67F2C9CF4EDB763F434B71DDDF6F53932EB6C662F0A779A99678E15E6ED7D4F3B4B282D973D4B0AD973442571EEC953EBC4505C9;
localparam G9_6 = 1024'h8869A86150E096B6565A3C70CC424AA50D897144B54A486337C49498C7622A3A8E756E60EE50A883919BA6CE2B81D6E4088B6B506AD7BFAA6EBC487D90C01FF96A0E6E16D6B855012A7F739B5C966AAB7BE4890291EBE105440B92764F9C3DA105688938966ACA5C10D7AB5EC2F9C4FE7FAA4443CE1623253D66A682CC6CFFEC;
localparam G9_7 = 1024'hE903248ECEA35C0175DD1674C42C2F4BCD1BC9FA89070DBFFD0A694C222D3D8EFEA0AE022FD63C82051F09B097BC52FECF86B095CA8C5ECB28E0857DC228151E8149923B8BD6BB5AAE5D087FB2EFD71998ECB76E94FE0DCC98C8A13C240B35AE158EB1126B54D02D845DDC1743B0D8E7BA14DC5D1D2D35D1EF139ED8446674AF;
localparam G9_8 = 1024'hD2834234E51165EE5C4EF15517D5528509EDDF99DDF712D21F1C3868769A2638051F169E27EDDBD94CFA85DF87CD6AB742AB8D1B861B876577D572D26B962E92AD5F628BDBA7501F58411BE04E5710C0B393CFB27BB049E8062072C1C9ED7BCE910B1365B65C005DD5FA019E608024FD4A8C1A41D79E213E9E0618032EB7815E;
localparam G10_1 = 1024'hD0D5550C36433A78B8E73DEBA50BB6D70AFD1E0AD800C39FED7206E10AAE9E329247E465BE1F60C42FD05463000AF629D5379CBE869B1BF1D85EE26D74DAE1F230920E307AE7D7ADDF0E80FAA37C6E42AB58E1D335863ECD206507319237ABE7E53442649215C16B8B6A042BD05BC678A8967CDA41DCE29C8950BE29E52A30FA;
localparam G10_2 = 1024'h43BA4B93DC7C549BC2239F96BFF547452D8B4D7C9117084F9F070CD7839FCBC94F185A81E4BB6D1C93541E6D097287C0BD70BFC16090A60757067544D57FCF9F0C9E33AB2118DC576DFC946BECAC23B2D93E1D5B72175398823C4918F8916EAB056C4FD94ED45266470E1AA1084206BBE5D62554B2130E97CBF16E1DA3B075B5;
localparam G10_3 = 1024'hC7BF2CE02A04964129D529AC269C20E7024B386D85CBF81D0402393BD718B6B7189941FCC1EDC72BE280526B063454B772DCE65CBC2C3DC23A172D30E819FC947EE891B1F3F6EF6AAFC512495CC1156D8BE6AC029DC5D1D1D24B18328B49A2A24952CC51C8B6F45335428422D794593D76CDF6E8B2EA0F0B76E75DC9B444B9B4;
localparam G10_4 = 1024'h2EBC2C83F375D1A6F807463B522BE8A8598D73718197B20C175578951E9D0489E174C03203BAAE91AF30735C97FE2B6355EB6ED9E48B5C9F58F58EA74470EC1B9975103F83AF500F31C685670103ECA9236BDE1417BA1326F91E37357DFEA07938E70AA706C96E423A1FF11D674736A5824EEDBA95B227C20AE44F47FF1954C5;
localparam G10_5 = 1024'hAFB905389867098E6934AC214E117BB7D43E4F20CC51B75B1BE75D61DAF157E47A90CBE8DB7708BA8D60FF4576502D0448A5A783CA3D402539CE191636AB7988FEC79B478D84C7979A5171CA6D27AB373EDED9C07503BCAC0DB85BB2D4D15B61FDF689E325915B5820A794709F393DB82F0FB519F20961C3E0869BD712BC3F1B;
localparam G10_6 = 1024'hEF2F24E09813BE117879F9BF30F55A03F93FF9F56DF438EC3CC8095361351BD32444DD557A4F6CDAB996FFA17AB99EFA6A98ECA05F245AD599BBFA08D86D63F737BBD947A4D89D52A0EE94E066EBAA0DD790826196FCDA3A3E2A3396067F019152111418F9103E4408DA8E1B425B825B70E6714DCD39F6AF1370C14450873305;
localparam G10_7 = 1024'hF87B3FF1DD2D2824DF10E38E82B324CB9500333D58A79CBEAB0902BD1EF2F5B4F9BC67E82CD0BF87846C6FA2AFE623BD5F826C2E5086AA66711B5D319F618F37E72F397323A163D5EDF3AF3FAFB135C0A8951F5FE4F85FE3F9B686FC762A461DB5332869D60766A5EBFC7714D4A015E053E066E6BC792188E6A962494E78C713;
localparam G10_8 = 1024'h22414395F088512D0F071297C3BF1F72DCB273D6C50BB3A2BB68DA5ABB6D994F1A8A1A5F16EB23D2C86D443DDB7F10CC4FCD4E05434C057D86CDAF8D5BA5F495AE16D560C9B71D1B639E78B5E993DAA84D6B900323BB28912B2AAC70CE42F18D7200B0FD53FCDE301F3682AFF6DA037827CE2F6ADFA8D058B4C081C838BA1CD8;
localparam G11_1 = 1024'hC5B00F91647A6720B71AFA0045CEB6A2C640D8B651DAECC3CB1662978E182FE2DECECD4EA4B7E9CB84CC72685BFBF45ACDBDA8CDD2E2997CADDC9E30BE52BB4C0D64D73147C9FC5B48381903D1B70F9A7485145E31A46C4CB00EA5E448691313EB5151C32626B956922BA2F6B4071360CBEBC960E64BD21E96CD25C409ED527E;
localparam G11_2 = 1024'h73E1AA4CA26BA8B49A96F56C8ECABBD9EA801F06E3CCCF2D55817340D7B0E43FD0E88FFB71D5BABBD4B6CC562150A85DD8D307371B66371FC30CB5BAAAD7A4800FC0CB6AB6805591D97BA4C6BD81CF5B0DDC699833DD90B26615B7560B4D7E1D26B54AD646860CBC045FF50BF6AAA815DE2746856EA74E33FD1E12D566A64C3E;
localparam G11_3 = 1024'hC71371AC71AF4D21DC1F73FA14E4AC642B6E3CDEDCF2FCC3DC86A05A41A9974EEBF597C4B82AAE2BFB0EB5DC1139AAE5CE639D9C10026C9FED5FA8D2064DA50BF689E63CE605A442457AFBA040912EC6B0AE1D7A83F82D0D71E62D36E2537FD21C1DF870792F8754872896C2D313947138B1344C33D874C4C0B08D20AF2D579E;
localparam G11_4 = 1024'h61D210EA2C3E77F4189EF580A123E41A76E124F86DE84CC81ED3AC638CB15DDB33D1DE7A6818B58D349CC2E60621175FB60371800EB18EB06C4005CDA0414795FE8B0FADC6B9BA279C707B9C5301255499786DC0C34E6397B7AA9193A302A50FEE60C4018F3054F9B1E795E72EE1ABD03132A684C741349E36FD96058BA02EB6;
localparam G11_5 = 1024'hD288899890EDAB3C7BF4950DA50899E6DB8D26FB51D3C58828A672DC9882C59D65243D2CED2083E5ED70D01562DD3FE317F1AF30483A6F188FA44A24AB479649145F77E4456005BC2FC50724A895C28822D9A1022B26D9357AD9416B8A8CF3C63937923B3886D80F0D115D1173835656A21F4E9878ABF203266D104C53FEC6E8;
localparam G11_6 = 1024'h3C979CAF0D253B90B2DC9AB895A50862DCCA2C3D3B9108FE89231CA0BFC78FD694F0D4BE64AB4BFB2CD446CF4C632E2383F7F529A6ECEBC02CE84D1367FEC91284EE2DD48EEAAFB7436EAE6432F0D9B608A24E8D11A59D5D4556E8FEDC9C54DD8F77F1DEBFF0062BF731CBDC1445387BFFF913FD5347DDD6299D8273D872702A;
localparam G11_7 = 1024'h2342B4846C21730E4F26362B722B0A4ED0D41BBB98D4A5B125C978E65133E0E879332632CDADCA05354B0339BC6FDE58182F12AC1F1C69FC425101C6E7AB009857EEDD1EEF2E74FC5743D768E75C5DA4BA8F1CD6F556EBDA4393EFB815DCF8F02C5B54CD33CD495C5B69D56B97F243CBC42F239BA44EA65891DA7C6626790BB0;
localparam G11_8 = 1024'hA55C3CAA65D282AFA7D06A86890B4A53ADEDC4492B15A839B8976B194BC331166AB0F4D06B9FE814C6B7239B8281EA7F07DCC96CE912140E2667A6CA29C25A52037E3BDC06670F23F73B50679EE61F67A253D28B661A0F6809DD001259EED99CFD81B9C824C1418DB0940ED4F88170AB20D4D4BB2F92A951849190E402724AA0;
localparam G12_1 = 1024'h204FD76BC8AB3CF4465263E30C01EA5E114BD548910135C58943A53A20E2D826218F99F8E75CBEB1610F141D9031869C6D8E54145405C3594DA2412A944D37D2C125086BECEED7E921E424BA8E8E0917A39C28966A1B72B57BBE26D1597648A9336A159738DD2A5E37B26C226C586948274796481A16DF23DE1C7FC931EDD219;
localparam G12_2 = 1024'h1B6DE14CA927E806ED3F401776863A728DEB7E05E202F37B526A661A7EABDB6C841DF0802E8AACACCDC56C2B272D29FF84FE8EC105E59691936EA829DEA6BBF32B4A164D960BA7FE6FCB8F24FAEFBEB42943838FC23427E92FC7AF990779727AA4FA48A7584897D521F584923512D38408E8562F5903BDE1C526794EBC3767A4;
localparam G12_3 = 1024'hA3AA71D6EFE407441E55C44F2329B170B9221078D3105763B8FA2C1EAF4F81617322F5E1CC31A5ADA6DC8428AD57CC62346D48B1124D20AD2084EE61A8FC4588C1893D38FB7CD310C26E1E2CA84A96AAF3EFAE1BCCBD69C8908BA14E071AFA50AA15CA830B67610449EE582AE6C147D86DFFB25BBF37350C3C3B9E66941D178C;
localparam G12_4 = 1024'hA46A27E3DBA91DA1B8BF4E26CB7A224D7EE3D80BB85B78B5408FA6FF3329D19B7CF6BE569708F1290FC338FA79E316DA09EB8FCEE7731A72452F79CC0CD68E9762DC07593766CC0EC1980BBA195F8D9D286E416220895DFCA5A3B8F6B828BA7CC1F6C39179F13972AA463C4F765F6D55F1A161E6717595D29C96AB487E27F413;
localparam G12_5 = 1024'h00795D64F8925631E1D67D9C20EE37ECBFE44BED04679AB4768CF38B7ED0EB480B13550387F7B9C369E643BB6F30048CF3E16D81A62DB6E6A7BE1EBC2A9EE8F9AB805D8709BEC88037796A51DB2D4FA3DA161DB43582EF21285BF19C539875A778A8681017F020E10B2114EBBF1B25121BCCF0FDA7505CE261C8297961E6CBE5;
localparam G12_6 = 1024'hEF94E9C253BA99C4522F1F46F60345E21DF4E42275569419AFA52B568169C2EA893B2ABB226A58A4564B2E51758D0D8A53443E8BBBF410DB00DCDA75C5E2D7B43D3E635A00CF241B90AE696B15F2FC3692CDFC9988EE4FBED43087658089E55946D559F2FCB5E122EAC6968033CC1CDB81E732001402BBC4EA1F0C6CC0D47A78;
localparam G12_7 = 1024'hF5B24A6FFAD18ACC2562433A59812281E7BC65DD36AEE6E84ABA791B74BCD479D1432219AFC683690CE2BA47B49DF331282AB07FBDE790E5FB4A292D15D0EB416059548D0762DBADC2F3962F98960AA5C4577A64A2416C0823A0C1D18792C7FE830D5CB977C7176C85B987A796FA46858EB1300BE729EC5F73785D94739E0ADA;
localparam G12_8 = 1024'h9308B6730E46C3EB90CBED7CB91046A680CEA38ECFF76B151132CDE7B9F6C5C12D64B83B4EECC4032FE959523D502366BF2823C96E0C8C8E1D8BFCB773E47AD7444AA0DCFE00F28B050D590A9D818A85CB10FED9E1A41C4BC64136D10D2F53C61CAE250767D8D78914BCB954B549A85BBEBD56BB697C1945BFF9C6DC8121A87A;
localparam G13_1 = 1024'hDFF8784B26817CAC72ABB22DF9E774072883EEDD803A82AA8FBB9142DC22CBDD108B8D24130838C8E84E0B981F281F79AEBC7C8E642B4ABBBC9735954ACF5125AAB49050AA07813C26F5F471E09DC1680E17C4EEF6C28E17696FF68AFCDB7DEF5B8272E0249AFA84CDF71E496B3EF87F12F8AFB227D8B1B5014D706C30C0CBBD;
localparam G13_2 = 1024'hA270CADD1BC31294A9FCEA16B528477588DBF86780D27C57573DBB901FF39DCB0029F94A8155588E18EC78BCD275BB5C3C16FE3BD284F53459917438060FBD7F0B9ECE57161AFB67A726EF73DE98A7AAFD9BEAC5AFD2249DEBF608D4FD02072522A15387C04955479817E2E2AEBB80E28719624DDF5F7A4E3FC34EDD2E53569C;
localparam G13_3 = 1024'h10E63EE5C13DAF5C157AE3927C0BEE26CB0D3D09764047453967975CE6C502CBBF95173D1B0A885AEDD502FEE067A8E60A4C094ECBBF363F2841AF59E3F9DB0A8C147831349C1961943FD2619368A6C5C44CB1F1F4B06963694FFD9D6360B2B73851EBE137CA8C06C44EDBE125961657441444A2167879656B2DF1B18568CC3C;
localparam G13_4 = 1024'h5A85E875862437E14CEF4C3CD7C15CF06C7C2A9820BBBB23FE081B8091BD24BCFD44BB8AAD56DCD04595146B5116E24514CE8EAC8D7E31C69A38F2665F54591CFC242D19570665A36F5BF4B91B2BB0D7F8AD1549F93E748D8807BFFD31531827E04E4F5FFFD3D739CCDA04E911D9DBC35F3BDA4DC4EA799DA65AF945A5EC9F6F;
localparam G13_5 = 1024'h3A4DE078CBB2328A82ECBB732AAFB17410CF23BD644E256720511CECD60BE50CDF7F46E66838B53B4C1BB251162152C290F28EA1D21A608CF7A51CEDD3AC4F75FDFB8945B2E9255137810021BB682D83BE768B24877162F3D9E956607149C26AD0C218B83DACF488A7EB0386348D5397EF2B28B4129C5CC10166C64E899319D4;
localparam G13_6 = 1024'h3193E8D954FE4993931A6BD38540150011189277351F0998F4990FD204C7C341B37C82B2C7F3ED8101D836B613657D0623812C4FC0092CDC00763132AF0797CD62231D4E406D2683D77151A22241A6628C7B6560D67EE5605DB2D79FB83A35926CEC3815F7938ECE0A8A06B9530767BEE2DE2B74336B3DFE510F3438EFF713DF;
localparam G13_7 = 1024'h106DC6B0A9F87575F55FB179648400657C33253FC56882CED5ECCE2D71692C45E43EC3478D2402D146B6D455719489468C49D9581D2E07D53910A7B21E9C483A82F9A7112FB28CBF7E4D1B77FB7BFED17E8EAE9A6FA71F1FE559DB4734D00B85B6D2A0E462BB31EA980EB7146830D26524CE148CE341B732B1E79964D8224BCC;
localparam G13_8 = 1024'h51F2DF994E8753BCF59FEAA2B4E9F1CA987F391EABF3F23D8388F36C4F7BA76347E47B31CE534C243A295A6CA12AFBE8F2BCC05C6BD334999F26439E7BE0E44736728CBBA762684613D6F70AA4751194138070B307513E6997597CBB2ACBDF98E17113A7AB28E917A62F69557A43C943ED0AF83F3EBBCF53AA070F55882FFE33;
localparam G14_1 = 1024'hD2C62B622393EBD7B9D62B5C46DCDB23D68E6B17D317415E3C7D0CA42D95426E6002A5C58BA0257DDC473BB780F4AE8389BF2FC1A3C41B80F8C267A424C99D02896182BE3D2CAE19480321A727F3C6C5C7DAD178FF971C1AFEA468023160391D460E79CED0D6B6F1EA9EBFFCDEF7EB69CFF6827C1C75106A6BF2F3F9C4B6EFD9;
localparam G14_2 = 1024'h95053BD28BA91952041D187937D509FF97F89DFFEC8ECB4B3DF53CBE3898675F47B019BCF053F4F62022383134BEEAEECED5EB14608ECD1A487050498CC60E9EB69C13259C9356F8DEE8D2283BE4278CE1F0D1414F2D9A48CDD74C23C8856D362B0ED42D9BFE6B99D4D64560770ECA843A016E2A2825091698D118ADD50DFBD4;
localparam G14_3 = 1024'h4BC27A27CFDCA686A7A4CB40D85A7D6627404DD151D88F6B6C6D1B0488B106F555DCE68361EDE8A4E3F0ECB137134485F8E52D3350CE392AEF4A46E18C52D05EACB3AB151EB7BAAFC997F6DBACF4967F9CBDC4B8C95DA0D242F5FB7B3C43B41F2E43ECBBF827B0C2084C854E917DB765A7634EB8C535DA40B27DE580FE432197;
localparam G14_4 = 1024'h25CA9FCACBA1C25430B44DC53C5D10670FEDBB82BF5D1DD0B9CAFDA75CD6CCFBE488768E264BE68EADFB8D62BEEB0E94E5B20ED59C562E0BE4C3C62B8F0A97272EBE05AF072BCF3C696FBEEBB05FD7E463F5F0761549718FCE0BADA5535BBB09976D162E201B49C27D97212840FDB81E0F31D5B2D6D6A86D30C392152CEC6B78;
localparam G14_5 = 1024'h7FA9E20561F5D35EAF105ED82B88D54A0172E85F0353912A7BB6CE512C31BDFA4FECE9737ECD84F0B396752654FE1CD5099D79DA62B45F7ED49D10DD0D0E6CFB0985A0D737BD7589FCE70E3B618FF7A089F4E11ED4AD7EE85AE214C3E2389C34EE0ED9BEB419B7752A57A484E31CF1A9CEDC94145FF08871E94D1C04FEFD3ACF;
localparam G14_6 = 1024'h2B5AD79A184B24557DD8DA5C10DFEA844E96CAF95750B971DF3B297C54B5AF3C4A7C26386F7B894796528C13DD5C48841C8840EC113945CE8C87FE83F404DA370E055D279AC035EFB7B1CBBDDCD4208761392DFA0EEBE30B302E70398C30F67107FF1BE35BEDBF3F9F898694589644BE683288FE039FDB83F01E75273C6ECC30;
localparam G14_7 = 1024'h763175618C7BD1349A5D0A5A0DC30D64B82A60F3EDDF0DC325FD7F6D13E0EAFAF94CE71BE8BEECD650A6E34764A3554C034426405001FC1309DC09CE16D4E153F05669FBC00E6E259568307411C2943BF2BEF7EC7D47131E685F601917CD990015468ED3DDA7841CEE625CA91BDACCB971E196AC4BD47CF813934390943D3386;
localparam G14_8 = 1024'h848BCE260584A605CBC1FFF1C05A67937D8765A654DF14A99EA78D5D2971CB245B2D704AC2C2CDE0862DD920EC37CCD16FBA2B681531E1A3CD12973A4E9D17FD47CC16138A34C0FD59383257A2B7E5185312668767E7EDE32C48DD050613040CAB7B632D29833A582D49677EDC99469704A813714C6E8729E59E2752A366BCCA;
localparam G15_1 = 1024'h33BDEA47E206055F05FCFA2ED7C7D66479A9798A9E8492B0EEB4CB138169B820DDC767D0EF3C908855153CB93E523524ADA80A327DDB04BC07F99DBE385F1BBE2ACF98E3BC2426E54F012197107D4347CC4B9737243E45D145B28A6B264BD91B513088D98832EEF3921C92A09A058F74E7944DE2FE93A54D4D65377AE5590C01;
localparam G15_2 = 1024'h90AC98B413A9D125A5E3DA85D23D29B1E37522FEE7C0F630BBF9DD6555749ADE8B47C989B46FB773D8C62A6C1B2A79FC3D04755C186D38A0F2A9D5500850AFA1B4B8B90F6CB84F76074EAF161B44C168D9513D0D9E252DB1AE7EBFB30A4FEA7F9B66FACE3252BC5A1819904FF1573A15B346EF7D917DDF19E8C264AFB040CB26;
localparam G15_3 = 1024'h57536A48937F6885084C0461411178720751A0FC5C54DC9010C7B475E666CC7113F7106B22B152998BBE75867940328E7359AE44AA07E257D4739696F99F49064A9697CB449C215B69EAE7DADBC50B63651FC5E473652CF6DC4475DAAAEBC1860FADF53AD2E49AC96523673201354381830AC85E043E892BEDFC418A1C77602A;
localparam G15_4 = 1024'h99EAD3855B0DE739CC04FDCCF4CB4467E5423EEB2D9AE1A4777D0E2EF5D7EE96C1A2DC2F7ED33B533D9356D97077A5AD78F669BC232E7216D1EDC2E34C2C5FE424A097A1E4B48AEEE9A058995EB6D73CBABC78C478333524DAFEE7E3E4D0D2E8EA266320481B98C4E602E76524E221E96233650754225288321EA0802FFB70ED;
localparam G15_5 = 1024'h2C0B29476A0EBC43B3CE4C8A907EF6EA574221EBF2BAC546D227B27CB753713C26C1FF3C3D8FCDC5F6797F629CF058540AE1B9F9D54DDFDCCC83A027940F5BB91641FD4D273BBDFFC25CCD6F9B5A9B1AB858B8F765D9B1CCF035AC0A6A6738F0DF5B51D754E1FB0AC172FFD22C748FD6DC9BB724B7DA5D6498151030A98818D0;
localparam G15_6 = 1024'h97BDF99DD76108CE8380887215423FD5A4FF664C76D69C159CC7F5194DCAE8EECDE5F1EC657EED929225BDA51349CBDA21C12F018A5C6AD0DAA27DB1D5AB0E5E31CB4A59E35137AD44BC6178E04775AC4C258C80CDAFFA401F081E5200145654112DB3FD7A5F07250DB1A99F967BBC25E121EF6A5F9C5B71E2D4512D85A08B00;
localparam G15_7 = 1024'h06FBF2CD7724DFC29DD352EAF6D34186ACABB8BF5DFA11CD033BC1C4187A6F9E14FCEA44958D50EAB84DD09F30D81E84BA3B48E93C578147DE97F4972AAE93EE21C5DBE8BB3ADDE6E0EA6AE8DE2D8EBAE603E04B26C2178C83B14C0BBFDEA3513905A8DF130F294070222F3E2AE8E48266847C90B1E1AE330B23714FE163C5BB;
localparam G15_8 = 1024'h2CBE168FF6803E943BB9B80603F5B752A3A91C5A437CEC621C79CC28F1D9776A24393948FA26DF81CBFAD60E0CC2FC8506124A636B6B3EB53AEFBE7AA0924956B2629B9C68B666D70C7DF94960E5A338E601AA6723037AF6742A37824E1D1C414938775E43C113997AD3CE79BE439351D16DB463A37CE82694DEF56FFCED14FF;
localparam G16_1 = 1024'h3426DFDB283B36981D8B3246ACC5D54976D19056833B23EE78F28B6AAE7B6E7E9ED558842F78BE2DD75B327394CB7B7AD6A421F30172830961D51B423E235813C422088BF996EB117447737B4C71C83CD4DAC20CB9F2AF53FF87F5656BD200EC6C7D80B47471A8E7CBBAFF0E0E5C052CEA1ABA4356E27E664CE1FBBA44B2CA6B;
localparam G16_2 = 1024'hDBDECE7442DC451EB8ECE8E5B00E0E2F0846D94951FC4E40490B7C377EBE93AA01E35547206DF3A9B77FAD82B7071DDE93B2798D1778B991257E93AB166F65831218ECF6968813F32147537F9EF347D1B8B15C24261D416351CD159664B2B5D1E982578B513166E0696ACEC0043503FF4752333618F6CC34BC621A7E09EBA5A1;
localparam G16_3 = 1024'h41216E0FC4E74D960EB9A288668F1F0249917A21FDBD34C9BD5034A5DA8C28DDC87DE14248720311E845396683A030930BC1CD89E0A5A2862B8BE3DC81A8B75C3845F2AE2E551C96CCCDCFF9FDBC3624EAFEF80018DFBFDF6673C99728AF2DCD78BA89CC5EB03FA57FA7E1896C9D43E6C9E6827FA77565270182AF4D43D3101D;
localparam G16_4 = 1024'hFD9695619F13D6848ACC26F3130F000ECB651CEB711630290692E45D125F48C9A222E323368339BA8CFBAFE54EA67D6FDE125D7B413266AF2808AA35D74093D04E2EBAFB0465990E82F1BF026D746EDD4501549EBF58697B1967EACF0A178E4F0D3104FD31758B617F44C5181ACD74946F1E0B02779065504F7A06792515FE3B;
localparam G16_5 = 1024'hFB7B506E8D172DBB893CC7AB8FC90997F640AF45A0C8F17BA9E21AF08F7FE673D2AA3D32A18083BBAB90AA05B943C1E0321B2BBDD9CD925CCE687B3DDD62A1D9C3FCAA422C363B3F2BF039C69EC273E74D0901AEFCFEB928E23F434DB9B88CFAED38A9748BEBFCF023020904566C26E31AF042710810AB75C8E47EA94463FF9E;
localparam G16_6 = 1024'h41E6250453E1FC44F93BF8A65BFFD0078CF6A65D4B8AD2F59632F4FA7F6D52284ED6E068FDB56C2B083A4AF81013FBFB5DC0BF286EB432A74F1D583F914143F1EE54CE5BED867C35721D0378B8E2C9C2069A4C9021395AE4861D88FAA0B6ECCB325A8E0106BA9FC7C4C195556EC8BFA54D470FF0B78D7EA8C6184286D3041A74;
localparam G16_7 = 1024'h41AA5D7FDAD019F22E5DDC3954B2038B08C0C5B3C77E48A2D3D8F49B4D64B50F622BB96698370CDD343E5C84FDC11236147BA5B5DDC91F0DAD621CF584D91354A43FAD039CF46E837B6921300B0015CEF6E409AE17969BDB0F5A53180B6D0FB9C7AB7E52A0A851C1D61943B73B3307BECC08A294753D8DBB6B7AAD74635C95E8;
localparam G16_8 = 1024'h1E46CDB452E52669E4321B73E4AE8FDF1EEA109819B398607AE3B4EC8A0EB63D7988B136679031A6D7C7152E18D4AB6D5368E9E08C961CC555E77666048AD1A60122D7556E9470AA45E83070090E20DEEA0DB44CFC037023A4FFCD546440F700CDE6016E35702C0CC5531BF9B8B6814C07E7B010EA3C00E8DFE3C17414BBAFCF;
/***********************************************************************************************************/
input clk;                             /*系统时钟*/
input rst_n;                           /*低电平异步复位信号*/

input [width-1:0] s_axis_tdata;        /*输入数据*/
input s_axis_tvalid;                   /*输入数据有效标志,高电平有效*/
output reg s_axis_tready;              /*向上游模块发送读请求或读确认信号,高电平有效*/

output reg [width-1:0] m_axis_tdata;   /*输出数据*/
output reg m_axis_tvalid;              /*输出数据有效标志,高电平有效*/
output reg m_axis_tlast;               /*码块结束标志位，每完成一个LDPC码块的输出拉高一次*/
input m_axis_tready;                   /*下游模块传来的读请求或读确认信号,高电平有效*/



/************************************************进行LDPC编码************************************************/
localparam STATE_waiting_valid=4'b1000;  /*等待valid信号*/
localparam STATE_data_out=4'b0100;       /*输出信息位*/
localparam STATE_waiting_ready=4'b0010;  /*等待ready信号*/
localparam STATE_check_out=4'b0001;      /*输出校验位*/

reg [3:0] state;               /*状态机*/
reg [$clog2(n):0] in_out_cnt;  /*输入/输出计数器*/
reg [n-k-1:0] g;               /*生成矩阵当前所在行*/
reg [n-k-1:0] check;           /*校验位*/
reg [width-1:0] s_tdata_reg;   /*输入寄存器*/
reg reg_flag;                  /*指示输入寄存器内是否有数据*/

wire [n-k-1:0] check_sub [width-1:0];
wire [n-k-1:0] check_reg;

assign check_sub[width-1]=m_axis_tdata[width-1]?g:0;
genvar i;
generate
for(i=0;i<=width-2;i=i+1)
begin
  assign check_sub[i]=m_axis_tdata[i]?({{g[sub_size*7+width-1-i-1:sub_size*7],g[sub_size*8-1:sub_size*7+width-1-i]},
                                        {g[sub_size*6+width-1-i-1:sub_size*6],g[sub_size*7-1:sub_size*6+width-1-i]},
                                        {g[sub_size*5+width-1-i-1:sub_size*5],g[sub_size*6-1:sub_size*5+width-1-i]},
                                        {g[sub_size*4+width-1-i-1:sub_size*4],g[sub_size*5-1:sub_size*4+width-1-i]},
                                        {g[sub_size*3+width-1-i-1:sub_size*3],g[sub_size*4-1:sub_size*3+width-1-i]},
                                        {g[sub_size*2+width-1-i-1:sub_size*2],g[sub_size*3-1:sub_size*2+width-1-i]},
                                        {g[sub_size*1+width-1-i-1:sub_size*1],g[sub_size*2-1:sub_size*1+width-1-i]},
                                        {g[sub_size*0+width-1-i-1:sub_size*0],g[sub_size*1-1:sub_size*0+width-1-i]}}):0;
end
endgenerate

generate
if(width==1)
  assign check_reg=check_sub[0];
else if(width==2)
  assign check_reg=check_sub[0]^check_sub[1];
else if(width==4)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3];
else if(width==8)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7];
else if(width==16)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15];
else if(width==32)
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15]^check_sub[16]^check_sub[17]^check_sub[18]^check_sub[19]^check_sub[20]^check_sub[21]^check_sub[22]^check_sub[23]^check_sub[24]^check_sub[25]^check_sub[26]^check_sub[27]^check_sub[28]^check_sub[29]^check_sub[30]^check_sub[31];
else
  assign check_reg=check_sub[0]^check_sub[1]^check_sub[2]^check_sub[3]^check_sub[4]^check_sub[5]^check_sub[6]^check_sub[7]^check_sub[8]^check_sub[9]^check_sub[10]^check_sub[11]^check_sub[12]^check_sub[13]^check_sub[14]^check_sub[15]^check_sub[16]^check_sub[17]^check_sub[18]^check_sub[19]^check_sub[20]^check_sub[21]^check_sub[22]^check_sub[23]^check_sub[24]^check_sub[25]^check_sub[26]^check_sub[27]^check_sub[28]^check_sub[29]^check_sub[30]^check_sub[31]^check_sub[32]^check_sub[33]^check_sub[34]^check_sub[35]^check_sub[36]^check_sub[37]^check_sub[38]^check_sub[39]^check_sub[40]^check_sub[41]^check_sub[42]^check_sub[43]^check_sub[44]^check_sub[45]^check_sub[46]^check_sub[47]^check_sub[48]^check_sub[49]^check_sub[50]^check_sub[51]^check_sub[52]^check_sub[53]^check_sub[54]^check_sub[55]^check_sub[56]^check_sub[57]^check_sub[58]^check_sub[59]^check_sub[60]^check_sub[61]^check_sub[62]^check_sub[63];
endgenerate

always@(posedge clk or negedge rst_n)
begin
  if(!rst_n)
    begin
      in_out_cnt<=0;
      g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
      check<=0;
      s_axis_tready<=0;
      s_tdata_reg<=0;
      reg_flag<=0;
      m_axis_tdata<=0;
      m_axis_tvalid<=0;
      m_axis_tlast<=0;
      state<=STATE_waiting_valid;
    end
  else
    begin
      case(state)
        STATE_waiting_valid : begin
                                s_axis_tready<=1;
                                if(s_axis_tready&&s_axis_tvalid) /*等待valid信号输入*/
                                  begin
                                    m_axis_tdata<=s_axis_tdata;
                                    m_axis_tvalid<=1;
                                    state<=STATE_data_out;
                                  end
                              end

        STATE_data_out : begin
                           if(m_axis_tready&&m_axis_tvalid)
                             begin
                               check<=check^check_reg; /*计算校验位*/
                               if(in_out_cnt==k-width) /*本码块的信息位输出完成*/
                                 begin
                                   in_out_cnt<=0;
                                   s_axis_tready<=0;
                                   m_axis_tdata<=m_axis_tdata;
                                   m_axis_tvalid<=0;
                                   state<=STATE_check_out;
                                   if(s_axis_tready&&s_axis_tvalid) /*输出本次信息位后,需继续输出校验位;若输入端具备有效数据,则将有效数据寄存*/
                                     begin
                                       s_tdata_reg<=s_axis_tdata;
                                       reg_flag<=1;
                                     end
                                 end
                               else
                                 begin
                                   in_out_cnt<=in_out_cnt+width;
                                   if(s_axis_tready&&s_axis_tvalid) /*输出本次信息位后,若输入端具备有效数据,则将有效数据输出*/
                                     begin
                                       m_axis_tdata<=s_axis_tdata;
                                       m_axis_tvalid<=1;
                                       state<=STATE_data_out;
                                     end
                                   else
                                     begin
                                       m_axis_tdata<=m_axis_tdata;
                                       m_axis_tvalid<=0;
                                       state<=STATE_waiting_valid;
                                     end
                                 end
                               case(in_out_cnt)
                                 sub_size*1-width : g<={G2_1,G2_2,G2_3,G2_4,G2_5,G2_6,G2_7,G2_8};
                                 sub_size*2-width : g<={G3_1,G3_2,G3_3,G3_4,G3_5,G3_6,G3_7,G3_8};
                                 sub_size*3-width : g<={G4_1,G4_2,G4_3,G4_4,G4_5,G4_6,G4_7,G4_8};
                                 sub_size*4-width : g<={G5_1,G5_2,G5_3,G5_4,G5_5,G5_6,G5_7,G5_8};
                                 sub_size*5-width : g<={G6_1,G6_2,G6_3,G6_4,G6_5,G6_6,G6_7,G6_8};
                                 sub_size*6-width : g<={G7_1,G7_2,G7_3,G7_4,G7_5,G7_6,G7_7,G7_8};
                                 sub_size*7-width : g<={G8_1,G8_2,G8_3,G8_4,G8_5,G8_6,G8_7,G8_8};
                                 sub_size*8-width : g<={G9_1,G9_2,G9_3,G9_4,G9_5,G9_6,G9_7,G9_8};
                                 sub_size*9-width : g<={G10_1,G10_2,G10_3,G10_4,G10_5,G10_6,G10_7,G10_8};
                                 sub_size*10-width: g<={G11_1,G11_2,G11_3,G11_4,G11_5,G11_6,G11_7,G11_8};
                                 sub_size*11-width: g<={G12_1,G12_2,G12_3,G12_4,G12_5,G12_6,G12_7,G12_8};
                                 sub_size*12-width: g<={G13_1,G13_2,G13_3,G13_4,G13_5,G13_6,G13_7,G13_8};
                                 sub_size*13-width: g<={G14_1,G14_2,G14_3,G14_4,G14_5,G14_6,G14_7,G14_8};
                                 sub_size*14-width: g<={G15_1,G15_2,G15_3,G15_4,G15_5,G15_6,G15_7,G15_8};
                                 sub_size*15-width: g<={G16_1,G16_2,G16_3,G16_4,G16_5,G16_6,G16_7,G16_8};
                                 sub_size*16-width: g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                                 default : g<={{g[sub_size*7+width-1:sub_size*7],g[sub_size*8-1:sub_size*7+width]},
                                               {g[sub_size*6+width-1:sub_size*6],g[sub_size*7-1:sub_size*6+width]},
                                               {g[sub_size*5+width-1:sub_size*5],g[sub_size*6-1:sub_size*5+width]},
                                               {g[sub_size*4+width-1:sub_size*4],g[sub_size*5-1:sub_size*4+width]},
                                               {g[sub_size*3+width-1:sub_size*3],g[sub_size*4-1:sub_size*3+width]},
                                               {g[sub_size*2+width-1:sub_size*2],g[sub_size*3-1:sub_size*2+width]},
                                               {g[sub_size*1+width-1:sub_size*1],g[sub_size*2-1:sub_size*1+width]},
                                               {g[sub_size*0+width-1:sub_size*0],g[sub_size*1-1:sub_size*0+width]}
                                              };
                               endcase
                             end
                           else /*后级模块不能接受数据,本次信息位输出未被后级模块取走*/
                             begin
                               s_axis_tready<=0;
                               state<=STATE_waiting_ready;
                               if(s_axis_tready&&s_axis_tvalid) /*本次输出未被取走,即使输入端具备有效数据,也不能将其更新至输出,只能寄存*/
                                 begin
                                   s_tdata_reg<=s_axis_tdata;
                                   reg_flag<=1;
                                 end
                             end
                         end
      
        STATE_waiting_ready : begin
                                if(m_axis_tready&&m_axis_tvalid)
                                  begin
                                    check<=check^check_reg;
                                    if(in_out_cnt==k-width)
                                      begin
                                        in_out_cnt<=0;
                                        m_axis_tdata<=m_axis_tdata;
                                        m_axis_tvalid<=0;
                                        state<=STATE_check_out;
                                      end
                                    else
                                      begin
                                        in_out_cnt<=in_out_cnt+width;
                                        s_axis_tready<=1;
                                        if(reg_flag==0)
                                          begin
                                            m_axis_tdata<=m_axis_tdata;
                                            m_axis_tvalid<=0;
                                            state<=STATE_waiting_valid;
                                          end
                                        else
                                          begin
                                            reg_flag<=0;
                                            m_axis_tdata<=s_tdata_reg;
                                            m_axis_tvalid<=1;
                                            state<=STATE_data_out;
                                          end
                                      end
                                    case(in_out_cnt)
                                      sub_size*1-width : g<={G2_1,G2_2,G2_3,G2_4,G2_5,G2_6,G2_7,G2_8};
                                      sub_size*2-width : g<={G3_1,G3_2,G3_3,G3_4,G3_5,G3_6,G3_7,G3_8};
                                      sub_size*3-width : g<={G4_1,G4_2,G4_3,G4_4,G4_5,G4_6,G4_7,G4_8};
                                      sub_size*4-width : g<={G5_1,G5_2,G5_3,G5_4,G5_5,G5_6,G5_7,G5_8};
                                      sub_size*5-width : g<={G6_1,G6_2,G6_3,G6_4,G6_5,G6_6,G6_7,G6_8};
                                      sub_size*6-width : g<={G7_1,G7_2,G7_3,G7_4,G7_5,G7_6,G7_7,G7_8};
                                      sub_size*7-width : g<={G8_1,G8_2,G8_3,G8_4,G8_5,G8_6,G8_7,G8_8};
                                      sub_size*8-width : g<={G9_1,G9_2,G9_3,G9_4,G9_5,G9_6,G9_7,G9_8};
                                      sub_size*9-width : g<={G10_1,G10_2,G10_3,G10_4,G10_5,G10_6,G10_7,G10_8};
                                      sub_size*10-width: g<={G11_1,G11_2,G11_3,G11_4,G11_5,G11_6,G11_7,G11_8};
                                      sub_size*11-width: g<={G12_1,G12_2,G12_3,G12_4,G12_5,G12_6,G12_7,G12_8};
                                      sub_size*12-width: g<={G13_1,G13_2,G13_3,G13_4,G13_5,G13_6,G13_7,G13_8};
                                      sub_size*13-width: g<={G14_1,G14_2,G14_3,G14_4,G14_5,G14_6,G14_7,G14_8};
                                      sub_size*14-width: g<={G15_1,G15_2,G15_3,G15_4,G15_5,G15_6,G15_7,G15_8};
                                      sub_size*15-width: g<={G16_1,G16_2,G16_3,G16_4,G16_5,G16_6,G16_7,G16_8};
                                      sub_size*16-width: g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                                      default : g<={{g[sub_size*7+width-1:sub_size*7],g[sub_size*8-1:sub_size*7+width]},
                                                    {g[sub_size*6+width-1:sub_size*6],g[sub_size*7-1:sub_size*6+width]},
                                                    {g[sub_size*5+width-1:sub_size*5],g[sub_size*6-1:sub_size*5+width]},
                                                    {g[sub_size*4+width-1:sub_size*4],g[sub_size*5-1:sub_size*4+width]},
                                                    {g[sub_size*3+width-1:sub_size*3],g[sub_size*4-1:sub_size*3+width]},
                                                    {g[sub_size*2+width-1:sub_size*2],g[sub_size*3-1:sub_size*2+width]},
                                                    {g[sub_size*1+width-1:sub_size*1],g[sub_size*2-1:sub_size*1+width]},
                                                    {g[sub_size*0+width-1:sub_size*0],g[sub_size*1-1:sub_size*0+width]}
                                                   };
                                    endcase
                                  end
                              end

        STATE_check_out : begin
                            if(!m_axis_tvalid)
                              begin
                                in_out_cnt<=0;
                                m_axis_tdata<=check[n-k-1:n-k-width];
                                m_axis_tvalid<=1;
                              end
                            else if(m_axis_tready&&m_axis_tvalid)
                              begin
                                if(in_out_cnt==n-k-width)
                                  begin
                                    in_out_cnt<=0;
                                    check<=0;
                                    s_axis_tready<=1;
                                    m_axis_tlast<=0;
                                    if(reg_flag)
                                      begin
                                        m_axis_tdata<=s_tdata_reg;
                                        reg_flag<=0;
                                        state<=STATE_data_out;
                                      end
                                    else
                                      begin
                                        m_axis_tdata<=m_axis_tdata;
                                        m_axis_tvalid<=0;
                                        state<=STATE_waiting_valid;
                                      end
                                  end
                                else if(in_out_cnt==n-k-2*width)
                                  begin
                                    in_out_cnt<=in_out_cnt+width;
                                    m_axis_tdata<=check[(n-k-1-in_out_cnt-width*2+1) +: width];
                                    m_axis_tlast<=1;
                                  end
                                else
                                  begin
                                    in_out_cnt<=in_out_cnt+width;
                                    m_axis_tdata<=check[(n-k-1-in_out_cnt-width*2+1) +: width];
                                  end
                              end
                          end
                          
        default : begin
                    in_out_cnt<=0;
                    g<={G1_1,G1_2,G1_3,G1_4,G1_5,G1_6,G1_7,G1_8};
                    check<=0;
                    s_axis_tready<=0;
                    m_axis_tdata<=0;
                    m_axis_tvalid<=0;
                    m_axis_tlast<=0;
                    state<=STATE_waiting_valid;            
                  end
      endcase
    end
end
/***********************************************************************************************************/

endmodule